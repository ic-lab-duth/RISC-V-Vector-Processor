module mul_(
input logic[31:0] a,
input logic[31:0] b,
output logic[63:0] res);
	logic in_0_0;
	logic in_0_1;
	logic in_1_0;
	logic in_0_2;
	logic in_1_1;
	logic in_2_0;
	logic in_0_3;
	logic in_1_2;
	logic in_2_1;
	logic in_3_0;
	logic in_0_4;
	logic in_1_3;
	logic in_2_2;
	logic in_3_1;
	logic in_4_0;
	logic in_0_5;
	logic in_1_4;
	logic in_2_3;
	logic in_3_2;
	logic in_4_1;
	logic in_5_0;
	logic in_0_6;
	logic in_1_5;
	logic in_2_4;
	logic in_3_3;
	logic in_4_2;
	logic in_5_1;
	logic in_6_0;
	logic in_0_7;
	logic in_1_6;
	logic in_2_5;
	logic in_3_4;
	logic in_4_3;
	logic in_5_2;
	logic in_6_1;
	logic in_7_0;
	logic in_0_8;
	logic in_1_7;
	logic in_2_6;
	logic in_3_5;
	logic in_4_4;
	logic in_5_3;
	logic in_6_2;
	logic in_7_1;
	logic in_8_0;
	logic in_0_9;
	logic in_1_8;
	logic in_2_7;
	logic in_3_6;
	logic in_4_5;
	logic in_5_4;
	logic in_6_3;
	logic in_7_2;
	logic in_8_1;
	logic in_9_0;
	logic in_0_10;
	logic in_1_9;
	logic in_2_8;
	logic in_3_7;
	logic in_4_6;
	logic in_5_5;
	logic in_6_4;
	logic in_7_3;
	logic in_8_2;
	logic in_9_1;
	logic in_10_0;
	logic in_0_11;
	logic in_1_10;
	logic in_2_9;
	logic in_3_8;
	logic in_4_7;
	logic in_5_6;
	logic in_6_5;
	logic in_7_4;
	logic in_8_3;
	logic in_9_2;
	logic in_10_1;
	logic in_11_0;
	logic in_0_12;
	logic in_1_11;
	logic in_2_10;
	logic in_3_9;
	logic in_4_8;
	logic in_5_7;
	logic in_6_6;
	logic in_7_5;
	logic in_8_4;
	logic in_9_3;
	logic in_10_2;
	logic in_11_1;
	logic in_12_0;
	logic in_0_13;
	logic in_1_12;
	logic in_2_11;
	logic in_3_10;
	logic in_4_9;
	logic in_5_8;
	logic in_6_7;
	logic in_7_6;
	logic in_8_5;
	logic in_9_4;
	logic in_10_3;
	logic in_11_2;
	logic in_12_1;
	logic in_13_0;
	logic in_0_14;
	logic in_1_13;
	logic in_2_12;
	logic in_3_11;
	logic in_4_10;
	logic in_5_9;
	logic in_6_8;
	logic in_7_7;
	logic in_8_6;
	logic in_9_5;
	logic in_10_4;
	logic in_11_3;
	logic in_12_2;
	logic in_13_1;
	logic in_14_0;
	logic in_0_15;
	logic in_1_14;
	logic in_2_13;
	logic in_3_12;
	logic in_4_11;
	logic in_5_10;
	logic in_6_9;
	logic in_7_8;
	logic in_8_7;
	logic in_9_6;
	logic in_10_5;
	logic in_11_4;
	logic in_12_3;
	logic in_13_2;
	logic in_14_1;
	logic in_15_0;
	logic in_0_16;
	logic in_1_15;
	logic in_2_14;
	logic in_3_13;
	logic in_4_12;
	logic in_5_11;
	logic in_6_10;
	logic in_7_9;
	logic in_8_8;
	logic in_9_7;
	logic in_10_6;
	logic in_11_5;
	logic in_12_4;
	logic in_13_3;
	logic in_14_2;
	logic in_15_1;
	logic in_16_0;
	logic in_0_17;
	logic in_1_16;
	logic in_2_15;
	logic in_3_14;
	logic in_4_13;
	logic in_5_12;
	logic in_6_11;
	logic in_7_10;
	logic in_8_9;
	logic in_9_8;
	logic in_10_7;
	logic in_11_6;
	logic in_12_5;
	logic in_13_4;
	logic in_14_3;
	logic in_15_2;
	logic in_16_1;
	logic in_17_0;
	logic in_0_18;
	logic in_1_17;
	logic in_2_16;
	logic in_3_15;
	logic in_4_14;
	logic in_5_13;
	logic in_6_12;
	logic in_7_11;
	logic in_8_10;
	logic in_9_9;
	logic in_10_8;
	logic in_11_7;
	logic in_12_6;
	logic in_13_5;
	logic in_14_4;
	logic in_15_3;
	logic in_16_2;
	logic in_17_1;
	logic in_18_0;
	logic in_0_19;
	logic in_1_18;
	logic in_2_17;
	logic in_3_16;
	logic in_4_15;
	logic in_5_14;
	logic in_6_13;
	logic in_7_12;
	logic in_8_11;
	logic in_9_10;
	logic in_10_9;
	logic in_11_8;
	logic in_12_7;
	logic in_13_6;
	logic in_14_5;
	logic in_15_4;
	logic in_16_3;
	logic in_17_2;
	logic in_18_1;
	logic in_19_0;
	logic in_0_20;
	logic in_1_19;
	logic in_2_18;
	logic in_3_17;
	logic in_4_16;
	logic in_5_15;
	logic in_6_14;
	logic in_7_13;
	logic in_8_12;
	logic in_9_11;
	logic in_10_10;
	logic in_11_9;
	logic in_12_8;
	logic in_13_7;
	logic in_14_6;
	logic in_15_5;
	logic in_16_4;
	logic in_17_3;
	logic in_18_2;
	logic in_19_1;
	logic in_20_0;
	logic in_0_21;
	logic in_1_20;
	logic in_2_19;
	logic in_3_18;
	logic in_4_17;
	logic in_5_16;
	logic in_6_15;
	logic in_7_14;
	logic in_8_13;
	logic in_9_12;
	logic in_10_11;
	logic in_11_10;
	logic in_12_9;
	logic in_13_8;
	logic in_14_7;
	logic in_15_6;
	logic in_16_5;
	logic in_17_4;
	logic in_18_3;
	logic in_19_2;
	logic in_20_1;
	logic in_21_0;
	logic in_0_22;
	logic in_1_21;
	logic in_2_20;
	logic in_3_19;
	logic in_4_18;
	logic in_5_17;
	logic in_6_16;
	logic in_7_15;
	logic in_8_14;
	logic in_9_13;
	logic in_10_12;
	logic in_11_11;
	logic in_12_10;
	logic in_13_9;
	logic in_14_8;
	logic in_15_7;
	logic in_16_6;
	logic in_17_5;
	logic in_18_4;
	logic in_19_3;
	logic in_20_2;
	logic in_21_1;
	logic in_22_0;
	logic in_0_23;
	logic in_1_22;
	logic in_2_21;
	logic in_3_20;
	logic in_4_19;
	logic in_5_18;
	logic in_6_17;
	logic in_7_16;
	logic in_8_15;
	logic in_9_14;
	logic in_10_13;
	logic in_11_12;
	logic in_12_11;
	logic in_13_10;
	logic in_14_9;
	logic in_15_8;
	logic in_16_7;
	logic in_17_6;
	logic in_18_5;
	logic in_19_4;
	logic in_20_3;
	logic in_21_2;
	logic in_22_1;
	logic in_23_0;
	logic in_0_24;
	logic in_1_23;
	logic in_2_22;
	logic in_3_21;
	logic in_4_20;
	logic in_5_19;
	logic in_6_18;
	logic in_7_17;
	logic in_8_16;
	logic in_9_15;
	logic in_10_14;
	logic in_11_13;
	logic in_12_12;
	logic in_13_11;
	logic in_14_10;
	logic in_15_9;
	logic in_16_8;
	logic in_17_7;
	logic in_18_6;
	logic in_19_5;
	logic in_20_4;
	logic in_21_3;
	logic in_22_2;
	logic in_23_1;
	logic in_24_0;
	logic in_0_25;
	logic in_1_24;
	logic in_2_23;
	logic in_3_22;
	logic in_4_21;
	logic in_5_20;
	logic in_6_19;
	logic in_7_18;
	logic in_8_17;
	logic in_9_16;
	logic in_10_15;
	logic in_11_14;
	logic in_12_13;
	logic in_13_12;
	logic in_14_11;
	logic in_15_10;
	logic in_16_9;
	logic in_17_8;
	logic in_18_7;
	logic in_19_6;
	logic in_20_5;
	logic in_21_4;
	logic in_22_3;
	logic in_23_2;
	logic in_24_1;
	logic in_25_0;
	logic in_0_26;
	logic in_1_25;
	logic in_2_24;
	logic in_3_23;
	logic in_4_22;
	logic in_5_21;
	logic in_6_20;
	logic in_7_19;
	logic in_8_18;
	logic in_9_17;
	logic in_10_16;
	logic in_11_15;
	logic in_12_14;
	logic in_13_13;
	logic in_14_12;
	logic in_15_11;
	logic in_16_10;
	logic in_17_9;
	logic in_18_8;
	logic in_19_7;
	logic in_20_6;
	logic in_21_5;
	logic in_22_4;
	logic in_23_3;
	logic in_24_2;
	logic in_25_1;
	logic in_26_0;
	logic in_0_27;
	logic in_1_26;
	logic in_2_25;
	logic in_3_24;
	logic in_4_23;
	logic in_5_22;
	logic in_6_21;
	logic in_7_20;
	logic in_8_19;
	logic in_9_18;
	logic in_10_17;
	logic in_11_16;
	logic in_12_15;
	logic in_13_14;
	logic in_14_13;
	logic in_15_12;
	logic in_16_11;
	logic in_17_10;
	logic in_18_9;
	logic in_19_8;
	logic in_20_7;
	logic in_21_6;
	logic in_22_5;
	logic in_23_4;
	logic in_24_3;
	logic in_25_2;
	logic in_26_1;
	logic in_27_0;
	logic in_0_28;
	logic in_1_27;
	logic in_2_26;
	logic in_3_25;
	logic in_4_24;
	logic in_5_23;
	logic in_6_22;
	logic in_7_21;
	logic in_8_20;
	logic in_9_19;
	logic in_10_18;
	logic in_11_17;
	logic in_12_16;
	logic in_13_15;
	logic in_14_14;
	logic in_15_13;
	logic in_16_12;
	logic in_17_11;
	logic in_18_10;
	logic in_19_9;
	logic in_20_8;
	logic in_21_7;
	logic in_22_6;
	logic in_23_5;
	logic in_24_4;
	logic in_25_3;
	logic in_26_2;
	logic in_27_1;
	logic in_28_0;
	logic in_0_29;
	logic in_1_28;
	logic in_2_27;
	logic in_3_26;
	logic in_4_25;
	logic in_5_24;
	logic in_6_23;
	logic in_7_22;
	logic in_8_21;
	logic in_9_20;
	logic in_10_19;
	logic in_11_18;
	logic in_12_17;
	logic in_13_16;
	logic in_14_15;
	logic in_15_14;
	logic in_16_13;
	logic in_17_12;
	logic in_18_11;
	logic in_19_10;
	logic in_20_9;
	logic in_21_8;
	logic in_22_7;
	logic in_23_6;
	logic in_24_5;
	logic in_25_4;
	logic in_26_3;
	logic in_27_2;
	logic in_28_1;
	logic in_29_0;
	logic in_0_30;
	logic in_1_29;
	logic in_2_28;
	logic in_3_27;
	logic in_4_26;
	logic in_5_25;
	logic in_6_24;
	logic in_7_23;
	logic in_8_22;
	logic in_9_21;
	logic in_10_20;
	logic in_11_19;
	logic in_12_18;
	logic in_13_17;
	logic in_14_16;
	logic in_15_15;
	logic in_16_14;
	logic in_17_13;
	logic in_18_12;
	logic in_19_11;
	logic in_20_10;
	logic in_21_9;
	logic in_22_8;
	logic in_23_7;
	logic in_24_6;
	logic in_25_5;
	logic in_26_4;
	logic in_27_3;
	logic in_28_2;
	logic in_29_1;
	logic in_30_0;
	logic in_0_31;
	logic in_1_30;
	logic in_2_29;
	logic in_3_28;
	logic in_4_27;
	logic in_5_26;
	logic in_6_25;
	logic in_7_24;
	logic in_8_23;
	logic in_9_22;
	logic in_10_21;
	logic in_11_20;
	logic in_12_19;
	logic in_13_18;
	logic in_14_17;
	logic in_15_16;
	logic in_16_15;
	logic in_17_14;
	logic in_18_13;
	logic in_19_12;
	logic in_20_11;
	logic in_21_10;
	logic in_22_9;
	logic in_23_8;
	logic in_24_7;
	logic in_25_6;
	logic in_26_5;
	logic in_27_4;
	logic in_28_3;
	logic in_29_2;
	logic in_30_1;
	logic in_31_0;
	logic in_1_31;
	logic in_2_30;
	logic in_3_29;
	logic in_4_28;
	logic in_5_27;
	logic in_6_26;
	logic in_7_25;
	logic in_8_24;
	logic in_9_23;
	logic in_10_22;
	logic in_11_21;
	logic in_12_20;
	logic in_13_19;
	logic in_14_18;
	logic in_15_17;
	logic in_16_16;
	logic in_17_15;
	logic in_18_14;
	logic in_19_13;
	logic in_20_12;
	logic in_21_11;
	logic in_22_10;
	logic in_23_9;
	logic in_24_8;
	logic in_25_7;
	logic in_26_6;
	logic in_27_5;
	logic in_28_4;
	logic in_29_3;
	logic in_30_2;
	logic in_31_1;
	logic in_2_31;
	logic in_3_30;
	logic in_4_29;
	logic in_5_28;
	logic in_6_27;
	logic in_7_26;
	logic in_8_25;
	logic in_9_24;
	logic in_10_23;
	logic in_11_22;
	logic in_12_21;
	logic in_13_20;
	logic in_14_19;
	logic in_15_18;
	logic in_16_17;
	logic in_17_16;
	logic in_18_15;
	logic in_19_14;
	logic in_20_13;
	logic in_21_12;
	logic in_22_11;
	logic in_23_10;
	logic in_24_9;
	logic in_25_8;
	logic in_26_7;
	logic in_27_6;
	logic in_28_5;
	logic in_29_4;
	logic in_30_3;
	logic in_31_2;
	logic in_3_31;
	logic in_4_30;
	logic in_5_29;
	logic in_6_28;
	logic in_7_27;
	logic in_8_26;
	logic in_9_25;
	logic in_10_24;
	logic in_11_23;
	logic in_12_22;
	logic in_13_21;
	logic in_14_20;
	logic in_15_19;
	logic in_16_18;
	logic in_17_17;
	logic in_18_16;
	logic in_19_15;
	logic in_20_14;
	logic in_21_13;
	logic in_22_12;
	logic in_23_11;
	logic in_24_10;
	logic in_25_9;
	logic in_26_8;
	logic in_27_7;
	logic in_28_6;
	logic in_29_5;
	logic in_30_4;
	logic in_31_3;
	logic in_4_31;
	logic in_5_30;
	logic in_6_29;
	logic in_7_28;
	logic in_8_27;
	logic in_9_26;
	logic in_10_25;
	logic in_11_24;
	logic in_12_23;
	logic in_13_22;
	logic in_14_21;
	logic in_15_20;
	logic in_16_19;
	logic in_17_18;
	logic in_18_17;
	logic in_19_16;
	logic in_20_15;
	logic in_21_14;
	logic in_22_13;
	logic in_23_12;
	logic in_24_11;
	logic in_25_10;
	logic in_26_9;
	logic in_27_8;
	logic in_28_7;
	logic in_29_6;
	logic in_30_5;
	logic in_31_4;
	logic in_5_31;
	logic in_6_30;
	logic in_7_29;
	logic in_8_28;
	logic in_9_27;
	logic in_10_26;
	logic in_11_25;
	logic in_12_24;
	logic in_13_23;
	logic in_14_22;
	logic in_15_21;
	logic in_16_20;
	logic in_17_19;
	logic in_18_18;
	logic in_19_17;
	logic in_20_16;
	logic in_21_15;
	logic in_22_14;
	logic in_23_13;
	logic in_24_12;
	logic in_25_11;
	logic in_26_10;
	logic in_27_9;
	logic in_28_8;
	logic in_29_7;
	logic in_30_6;
	logic in_31_5;
	logic in_6_31;
	logic in_7_30;
	logic in_8_29;
	logic in_9_28;
	logic in_10_27;
	logic in_11_26;
	logic in_12_25;
	logic in_13_24;
	logic in_14_23;
	logic in_15_22;
	logic in_16_21;
	logic in_17_20;
	logic in_18_19;
	logic in_19_18;
	logic in_20_17;
	logic in_21_16;
	logic in_22_15;
	logic in_23_14;
	logic in_24_13;
	logic in_25_12;
	logic in_26_11;
	logic in_27_10;
	logic in_28_9;
	logic in_29_8;
	logic in_30_7;
	logic in_31_6;
	logic in_7_31;
	logic in_8_30;
	logic in_9_29;
	logic in_10_28;
	logic in_11_27;
	logic in_12_26;
	logic in_13_25;
	logic in_14_24;
	logic in_15_23;
	logic in_16_22;
	logic in_17_21;
	logic in_18_20;
	logic in_19_19;
	logic in_20_18;
	logic in_21_17;
	logic in_22_16;
	logic in_23_15;
	logic in_24_14;
	logic in_25_13;
	logic in_26_12;
	logic in_27_11;
	logic in_28_10;
	logic in_29_9;
	logic in_30_8;
	logic in_31_7;
	logic in_8_31;
	logic in_9_30;
	logic in_10_29;
	logic in_11_28;
	logic in_12_27;
	logic in_13_26;
	logic in_14_25;
	logic in_15_24;
	logic in_16_23;
	logic in_17_22;
	logic in_18_21;
	logic in_19_20;
	logic in_20_19;
	logic in_21_18;
	logic in_22_17;
	logic in_23_16;
	logic in_24_15;
	logic in_25_14;
	logic in_26_13;
	logic in_27_12;
	logic in_28_11;
	logic in_29_10;
	logic in_30_9;
	logic in_31_8;
	logic in_9_31;
	logic in_10_30;
	logic in_11_29;
	logic in_12_28;
	logic in_13_27;
	logic in_14_26;
	logic in_15_25;
	logic in_16_24;
	logic in_17_23;
	logic in_18_22;
	logic in_19_21;
	logic in_20_20;
	logic in_21_19;
	logic in_22_18;
	logic in_23_17;
	logic in_24_16;
	logic in_25_15;
	logic in_26_14;
	logic in_27_13;
	logic in_28_12;
	logic in_29_11;
	logic in_30_10;
	logic in_31_9;
	logic in_10_31;
	logic in_11_30;
	logic in_12_29;
	logic in_13_28;
	logic in_14_27;
	logic in_15_26;
	logic in_16_25;
	logic in_17_24;
	logic in_18_23;
	logic in_19_22;
	logic in_20_21;
	logic in_21_20;
	logic in_22_19;
	logic in_23_18;
	logic in_24_17;
	logic in_25_16;
	logic in_26_15;
	logic in_27_14;
	logic in_28_13;
	logic in_29_12;
	logic in_30_11;
	logic in_31_10;
	logic in_11_31;
	logic in_12_30;
	logic in_13_29;
	logic in_14_28;
	logic in_15_27;
	logic in_16_26;
	logic in_17_25;
	logic in_18_24;
	logic in_19_23;
	logic in_20_22;
	logic in_21_21;
	logic in_22_20;
	logic in_23_19;
	logic in_24_18;
	logic in_25_17;
	logic in_26_16;
	logic in_27_15;
	logic in_28_14;
	logic in_29_13;
	logic in_30_12;
	logic in_31_11;
	logic in_12_31;
	logic in_13_30;
	logic in_14_29;
	logic in_15_28;
	logic in_16_27;
	logic in_17_26;
	logic in_18_25;
	logic in_19_24;
	logic in_20_23;
	logic in_21_22;
	logic in_22_21;
	logic in_23_20;
	logic in_24_19;
	logic in_25_18;
	logic in_26_17;
	logic in_27_16;
	logic in_28_15;
	logic in_29_14;
	logic in_30_13;
	logic in_31_12;
	logic in_13_31;
	logic in_14_30;
	logic in_15_29;
	logic in_16_28;
	logic in_17_27;
	logic in_18_26;
	logic in_19_25;
	logic in_20_24;
	logic in_21_23;
	logic in_22_22;
	logic in_23_21;
	logic in_24_20;
	logic in_25_19;
	logic in_26_18;
	logic in_27_17;
	logic in_28_16;
	logic in_29_15;
	logic in_30_14;
	logic in_31_13;
	logic in_14_31;
	logic in_15_30;
	logic in_16_29;
	logic in_17_28;
	logic in_18_27;
	logic in_19_26;
	logic in_20_25;
	logic in_21_24;
	logic in_22_23;
	logic in_23_22;
	logic in_24_21;
	logic in_25_20;
	logic in_26_19;
	logic in_27_18;
	logic in_28_17;
	logic in_29_16;
	logic in_30_15;
	logic in_31_14;
	logic in_15_31;
	logic in_16_30;
	logic in_17_29;
	logic in_18_28;
	logic in_19_27;
	logic in_20_26;
	logic in_21_25;
	logic in_22_24;
	logic in_23_23;
	logic in_24_22;
	logic in_25_21;
	logic in_26_20;
	logic in_27_19;
	logic in_28_18;
	logic in_29_17;
	logic in_30_16;
	logic in_31_15;
	logic in_16_31;
	logic in_17_30;
	logic in_18_29;
	logic in_19_28;
	logic in_20_27;
	logic in_21_26;
	logic in_22_25;
	logic in_23_24;
	logic in_24_23;
	logic in_25_22;
	logic in_26_21;
	logic in_27_20;
	logic in_28_19;
	logic in_29_18;
	logic in_30_17;
	logic in_31_16;
	logic in_17_31;
	logic in_18_30;
	logic in_19_29;
	logic in_20_28;
	logic in_21_27;
	logic in_22_26;
	logic in_23_25;
	logic in_24_24;
	logic in_25_23;
	logic in_26_22;
	logic in_27_21;
	logic in_28_20;
	logic in_29_19;
	logic in_30_18;
	logic in_31_17;
	logic in_18_31;
	logic in_19_30;
	logic in_20_29;
	logic in_21_28;
	logic in_22_27;
	logic in_23_26;
	logic in_24_25;
	logic in_25_24;
	logic in_26_23;
	logic in_27_22;
	logic in_28_21;
	logic in_29_20;
	logic in_30_19;
	logic in_31_18;
	logic in_19_31;
	logic in_20_30;
	logic in_21_29;
	logic in_22_28;
	logic in_23_27;
	logic in_24_26;
	logic in_25_25;
	logic in_26_24;
	logic in_27_23;
	logic in_28_22;
	logic in_29_21;
	logic in_30_20;
	logic in_31_19;
	logic in_20_31;
	logic in_21_30;
	logic in_22_29;
	logic in_23_28;
	logic in_24_27;
	logic in_25_26;
	logic in_26_25;
	logic in_27_24;
	logic in_28_23;
	logic in_29_22;
	logic in_30_21;
	logic in_31_20;
	logic in_21_31;
	logic in_22_30;
	logic in_23_29;
	logic in_24_28;
	logic in_25_27;
	logic in_26_26;
	logic in_27_25;
	logic in_28_24;
	logic in_29_23;
	logic in_30_22;
	logic in_31_21;
	logic in_22_31;
	logic in_23_30;
	logic in_24_29;
	logic in_25_28;
	logic in_26_27;
	logic in_27_26;
	logic in_28_25;
	logic in_29_24;
	logic in_30_23;
	logic in_31_22;
	logic in_23_31;
	logic in_24_30;
	logic in_25_29;
	logic in_26_28;
	logic in_27_27;
	logic in_28_26;
	logic in_29_25;
	logic in_30_24;
	logic in_31_23;
	logic in_24_31;
	logic in_25_30;
	logic in_26_29;
	logic in_27_28;
	logic in_28_27;
	logic in_29_26;
	logic in_30_25;
	logic in_31_24;
	logic in_25_31;
	logic in_26_30;
	logic in_27_29;
	logic in_28_28;
	logic in_29_27;
	logic in_30_26;
	logic in_31_25;
	logic in_26_31;
	logic in_27_30;
	logic in_28_29;
	logic in_29_28;
	logic in_30_27;
	logic in_31_26;
	logic in_27_31;
	logic in_28_30;
	logic in_29_29;
	logic in_30_28;
	logic in_31_27;
	logic in_28_31;
	logic in_29_30;
	logic in_30_29;
	logic in_31_28;
	logic in_29_31;
	logic in_30_30;
	logic in_31_29;
	logic in_30_31;
	logic in_31_30;
	logic in_31_31;

	assign in_0_0 = a[0]&b[0];
	assign in_1_0 = a[1]&b[0];
	assign in_2_0 = a[2]&b[0];
	assign in_3_0 = a[3]&b[0];
	assign in_4_0 = a[4]&b[0];
	assign in_5_0 = a[5]&b[0];
	assign in_6_0 = a[6]&b[0];
	assign in_7_0 = a[7]&b[0];
	assign in_8_0 = a[8]&b[0];
	assign in_9_0 = a[9]&b[0];
	assign in_10_0 = a[10]&b[0];
	assign in_11_0 = a[11]&b[0];
	assign in_12_0 = a[12]&b[0];
	assign in_13_0 = a[13]&b[0];
	assign in_14_0 = a[14]&b[0];
	assign in_15_0 = a[15]&b[0];
	assign in_16_0 = a[16]&b[0];
	assign in_17_0 = a[17]&b[0];
	assign in_18_0 = a[18]&b[0];
	assign in_19_0 = a[19]&b[0];
	assign in_20_0 = a[20]&b[0];
	assign in_21_0 = a[21]&b[0];
	assign in_22_0 = a[22]&b[0];
	assign in_23_0 = a[23]&b[0];
	assign in_24_0 = a[24]&b[0];
	assign in_25_0 = a[25]&b[0];
	assign in_26_0 = a[26]&b[0];
	assign in_27_0 = a[27]&b[0];
	assign in_28_0 = a[28]&b[0];
	assign in_29_0 = a[29]&b[0];
	assign in_30_0 = a[30]&b[0];
	assign in_31_0 = a[31]&b[0];
	assign in_0_1 = a[0]&b[1];
	assign in_1_1 = a[1]&b[1];
	assign in_2_1 = a[2]&b[1];
	assign in_3_1 = a[3]&b[1];
	assign in_4_1 = a[4]&b[1];
	assign in_5_1 = a[5]&b[1];
	assign in_6_1 = a[6]&b[1];
	assign in_7_1 = a[7]&b[1];
	assign in_8_1 = a[8]&b[1];
	assign in_9_1 = a[9]&b[1];
	assign in_10_1 = a[10]&b[1];
	assign in_11_1 = a[11]&b[1];
	assign in_12_1 = a[12]&b[1];
	assign in_13_1 = a[13]&b[1];
	assign in_14_1 = a[14]&b[1];
	assign in_15_1 = a[15]&b[1];
	assign in_16_1 = a[16]&b[1];
	assign in_17_1 = a[17]&b[1];
	assign in_18_1 = a[18]&b[1];
	assign in_19_1 = a[19]&b[1];
	assign in_20_1 = a[20]&b[1];
	assign in_21_1 = a[21]&b[1];
	assign in_22_1 = a[22]&b[1];
	assign in_23_1 = a[23]&b[1];
	assign in_24_1 = a[24]&b[1];
	assign in_25_1 = a[25]&b[1];
	assign in_26_1 = a[26]&b[1];
	assign in_27_1 = a[27]&b[1];
	assign in_28_1 = a[28]&b[1];
	assign in_29_1 = a[29]&b[1];
	assign in_30_1 = a[30]&b[1];
	assign in_31_1 = a[31]&b[1];
	assign in_0_2 = a[0]&b[2];
	assign in_1_2 = a[1]&b[2];
	assign in_2_2 = a[2]&b[2];
	assign in_3_2 = a[3]&b[2];
	assign in_4_2 = a[4]&b[2];
	assign in_5_2 = a[5]&b[2];
	assign in_6_2 = a[6]&b[2];
	assign in_7_2 = a[7]&b[2];
	assign in_8_2 = a[8]&b[2];
	assign in_9_2 = a[9]&b[2];
	assign in_10_2 = a[10]&b[2];
	assign in_11_2 = a[11]&b[2];
	assign in_12_2 = a[12]&b[2];
	assign in_13_2 = a[13]&b[2];
	assign in_14_2 = a[14]&b[2];
	assign in_15_2 = a[15]&b[2];
	assign in_16_2 = a[16]&b[2];
	assign in_17_2 = a[17]&b[2];
	assign in_18_2 = a[18]&b[2];
	assign in_19_2 = a[19]&b[2];
	assign in_20_2 = a[20]&b[2];
	assign in_21_2 = a[21]&b[2];
	assign in_22_2 = a[22]&b[2];
	assign in_23_2 = a[23]&b[2];
	assign in_24_2 = a[24]&b[2];
	assign in_25_2 = a[25]&b[2];
	assign in_26_2 = a[26]&b[2];
	assign in_27_2 = a[27]&b[2];
	assign in_28_2 = a[28]&b[2];
	assign in_29_2 = a[29]&b[2];
	assign in_30_2 = a[30]&b[2];
	assign in_31_2 = a[31]&b[2];
	assign in_0_3 = a[0]&b[3];
	assign in_1_3 = a[1]&b[3];
	assign in_2_3 = a[2]&b[3];
	assign in_3_3 = a[3]&b[3];
	assign in_4_3 = a[4]&b[3];
	assign in_5_3 = a[5]&b[3];
	assign in_6_3 = a[6]&b[3];
	assign in_7_3 = a[7]&b[3];
	assign in_8_3 = a[8]&b[3];
	assign in_9_3 = a[9]&b[3];
	assign in_10_3 = a[10]&b[3];
	assign in_11_3 = a[11]&b[3];
	assign in_12_3 = a[12]&b[3];
	assign in_13_3 = a[13]&b[3];
	assign in_14_3 = a[14]&b[3];
	assign in_15_3 = a[15]&b[3];
	assign in_16_3 = a[16]&b[3];
	assign in_17_3 = a[17]&b[3];
	assign in_18_3 = a[18]&b[3];
	assign in_19_3 = a[19]&b[3];
	assign in_20_3 = a[20]&b[3];
	assign in_21_3 = a[21]&b[3];
	assign in_22_3 = a[22]&b[3];
	assign in_23_3 = a[23]&b[3];
	assign in_24_3 = a[24]&b[3];
	assign in_25_3 = a[25]&b[3];
	assign in_26_3 = a[26]&b[3];
	assign in_27_3 = a[27]&b[3];
	assign in_28_3 = a[28]&b[3];
	assign in_29_3 = a[29]&b[3];
	assign in_30_3 = a[30]&b[3];
	assign in_31_3 = a[31]&b[3];
	assign in_0_4 = a[0]&b[4];
	assign in_1_4 = a[1]&b[4];
	assign in_2_4 = a[2]&b[4];
	assign in_3_4 = a[3]&b[4];
	assign in_4_4 = a[4]&b[4];
	assign in_5_4 = a[5]&b[4];
	assign in_6_4 = a[6]&b[4];
	assign in_7_4 = a[7]&b[4];
	assign in_8_4 = a[8]&b[4];
	assign in_9_4 = a[9]&b[4];
	assign in_10_4 = a[10]&b[4];
	assign in_11_4 = a[11]&b[4];
	assign in_12_4 = a[12]&b[4];
	assign in_13_4 = a[13]&b[4];
	assign in_14_4 = a[14]&b[4];
	assign in_15_4 = a[15]&b[4];
	assign in_16_4 = a[16]&b[4];
	assign in_17_4 = a[17]&b[4];
	assign in_18_4 = a[18]&b[4];
	assign in_19_4 = a[19]&b[4];
	assign in_20_4 = a[20]&b[4];
	assign in_21_4 = a[21]&b[4];
	assign in_22_4 = a[22]&b[4];
	assign in_23_4 = a[23]&b[4];
	assign in_24_4 = a[24]&b[4];
	assign in_25_4 = a[25]&b[4];
	assign in_26_4 = a[26]&b[4];
	assign in_27_4 = a[27]&b[4];
	assign in_28_4 = a[28]&b[4];
	assign in_29_4 = a[29]&b[4];
	assign in_30_4 = a[30]&b[4];
	assign in_31_4 = a[31]&b[4];
	assign in_0_5 = a[0]&b[5];
	assign in_1_5 = a[1]&b[5];
	assign in_2_5 = a[2]&b[5];
	assign in_3_5 = a[3]&b[5];
	assign in_4_5 = a[4]&b[5];
	assign in_5_5 = a[5]&b[5];
	assign in_6_5 = a[6]&b[5];
	assign in_7_5 = a[7]&b[5];
	assign in_8_5 = a[8]&b[5];
	assign in_9_5 = a[9]&b[5];
	assign in_10_5 = a[10]&b[5];
	assign in_11_5 = a[11]&b[5];
	assign in_12_5 = a[12]&b[5];
	assign in_13_5 = a[13]&b[5];
	assign in_14_5 = a[14]&b[5];
	assign in_15_5 = a[15]&b[5];
	assign in_16_5 = a[16]&b[5];
	assign in_17_5 = a[17]&b[5];
	assign in_18_5 = a[18]&b[5];
	assign in_19_5 = a[19]&b[5];
	assign in_20_5 = a[20]&b[5];
	assign in_21_5 = a[21]&b[5];
	assign in_22_5 = a[22]&b[5];
	assign in_23_5 = a[23]&b[5];
	assign in_24_5 = a[24]&b[5];
	assign in_25_5 = a[25]&b[5];
	assign in_26_5 = a[26]&b[5];
	assign in_27_5 = a[27]&b[5];
	assign in_28_5 = a[28]&b[5];
	assign in_29_5 = a[29]&b[5];
	assign in_30_5 = a[30]&b[5];
	assign in_31_5 = a[31]&b[5];
	assign in_0_6 = a[0]&b[6];
	assign in_1_6 = a[1]&b[6];
	assign in_2_6 = a[2]&b[6];
	assign in_3_6 = a[3]&b[6];
	assign in_4_6 = a[4]&b[6];
	assign in_5_6 = a[5]&b[6];
	assign in_6_6 = a[6]&b[6];
	assign in_7_6 = a[7]&b[6];
	assign in_8_6 = a[8]&b[6];
	assign in_9_6 = a[9]&b[6];
	assign in_10_6 = a[10]&b[6];
	assign in_11_6 = a[11]&b[6];
	assign in_12_6 = a[12]&b[6];
	assign in_13_6 = a[13]&b[6];
	assign in_14_6 = a[14]&b[6];
	assign in_15_6 = a[15]&b[6];
	assign in_16_6 = a[16]&b[6];
	assign in_17_6 = a[17]&b[6];
	assign in_18_6 = a[18]&b[6];
	assign in_19_6 = a[19]&b[6];
	assign in_20_6 = a[20]&b[6];
	assign in_21_6 = a[21]&b[6];
	assign in_22_6 = a[22]&b[6];
	assign in_23_6 = a[23]&b[6];
	assign in_24_6 = a[24]&b[6];
	assign in_25_6 = a[25]&b[6];
	assign in_26_6 = a[26]&b[6];
	assign in_27_6 = a[27]&b[6];
	assign in_28_6 = a[28]&b[6];
	assign in_29_6 = a[29]&b[6];
	assign in_30_6 = a[30]&b[6];
	assign in_31_6 = a[31]&b[6];
	assign in_0_7 = a[0]&b[7];
	assign in_1_7 = a[1]&b[7];
	assign in_2_7 = a[2]&b[7];
	assign in_3_7 = a[3]&b[7];
	assign in_4_7 = a[4]&b[7];
	assign in_5_7 = a[5]&b[7];
	assign in_6_7 = a[6]&b[7];
	assign in_7_7 = a[7]&b[7];
	assign in_8_7 = a[8]&b[7];
	assign in_9_7 = a[9]&b[7];
	assign in_10_7 = a[10]&b[7];
	assign in_11_7 = a[11]&b[7];
	assign in_12_7 = a[12]&b[7];
	assign in_13_7 = a[13]&b[7];
	assign in_14_7 = a[14]&b[7];
	assign in_15_7 = a[15]&b[7];
	assign in_16_7 = a[16]&b[7];
	assign in_17_7 = a[17]&b[7];
	assign in_18_7 = a[18]&b[7];
	assign in_19_7 = a[19]&b[7];
	assign in_20_7 = a[20]&b[7];
	assign in_21_7 = a[21]&b[7];
	assign in_22_7 = a[22]&b[7];
	assign in_23_7 = a[23]&b[7];
	assign in_24_7 = a[24]&b[7];
	assign in_25_7 = a[25]&b[7];
	assign in_26_7 = a[26]&b[7];
	assign in_27_7 = a[27]&b[7];
	assign in_28_7 = a[28]&b[7];
	assign in_29_7 = a[29]&b[7];
	assign in_30_7 = a[30]&b[7];
	assign in_31_7 = a[31]&b[7];
	assign in_0_8 = a[0]&b[8];
	assign in_1_8 = a[1]&b[8];
	assign in_2_8 = a[2]&b[8];
	assign in_3_8 = a[3]&b[8];
	assign in_4_8 = a[4]&b[8];
	assign in_5_8 = a[5]&b[8];
	assign in_6_8 = a[6]&b[8];
	assign in_7_8 = a[7]&b[8];
	assign in_8_8 = a[8]&b[8];
	assign in_9_8 = a[9]&b[8];
	assign in_10_8 = a[10]&b[8];
	assign in_11_8 = a[11]&b[8];
	assign in_12_8 = a[12]&b[8];
	assign in_13_8 = a[13]&b[8];
	assign in_14_8 = a[14]&b[8];
	assign in_15_8 = a[15]&b[8];
	assign in_16_8 = a[16]&b[8];
	assign in_17_8 = a[17]&b[8];
	assign in_18_8 = a[18]&b[8];
	assign in_19_8 = a[19]&b[8];
	assign in_20_8 = a[20]&b[8];
	assign in_21_8 = a[21]&b[8];
	assign in_22_8 = a[22]&b[8];
	assign in_23_8 = a[23]&b[8];
	assign in_24_8 = a[24]&b[8];
	assign in_25_8 = a[25]&b[8];
	assign in_26_8 = a[26]&b[8];
	assign in_27_8 = a[27]&b[8];
	assign in_28_8 = a[28]&b[8];
	assign in_29_8 = a[29]&b[8];
	assign in_30_8 = a[30]&b[8];
	assign in_31_8 = a[31]&b[8];
	assign in_0_9 = a[0]&b[9];
	assign in_1_9 = a[1]&b[9];
	assign in_2_9 = a[2]&b[9];
	assign in_3_9 = a[3]&b[9];
	assign in_4_9 = a[4]&b[9];
	assign in_5_9 = a[5]&b[9];
	assign in_6_9 = a[6]&b[9];
	assign in_7_9 = a[7]&b[9];
	assign in_8_9 = a[8]&b[9];
	assign in_9_9 = a[9]&b[9];
	assign in_10_9 = a[10]&b[9];
	assign in_11_9 = a[11]&b[9];
	assign in_12_9 = a[12]&b[9];
	assign in_13_9 = a[13]&b[9];
	assign in_14_9 = a[14]&b[9];
	assign in_15_9 = a[15]&b[9];
	assign in_16_9 = a[16]&b[9];
	assign in_17_9 = a[17]&b[9];
	assign in_18_9 = a[18]&b[9];
	assign in_19_9 = a[19]&b[9];
	assign in_20_9 = a[20]&b[9];
	assign in_21_9 = a[21]&b[9];
	assign in_22_9 = a[22]&b[9];
	assign in_23_9 = a[23]&b[9];
	assign in_24_9 = a[24]&b[9];
	assign in_25_9 = a[25]&b[9];
	assign in_26_9 = a[26]&b[9];
	assign in_27_9 = a[27]&b[9];
	assign in_28_9 = a[28]&b[9];
	assign in_29_9 = a[29]&b[9];
	assign in_30_9 = a[30]&b[9];
	assign in_31_9 = a[31]&b[9];
	assign in_0_10 = a[0]&b[10];
	assign in_1_10 = a[1]&b[10];
	assign in_2_10 = a[2]&b[10];
	assign in_3_10 = a[3]&b[10];
	assign in_4_10 = a[4]&b[10];
	assign in_5_10 = a[5]&b[10];
	assign in_6_10 = a[6]&b[10];
	assign in_7_10 = a[7]&b[10];
	assign in_8_10 = a[8]&b[10];
	assign in_9_10 = a[9]&b[10];
	assign in_10_10 = a[10]&b[10];
	assign in_11_10 = a[11]&b[10];
	assign in_12_10 = a[12]&b[10];
	assign in_13_10 = a[13]&b[10];
	assign in_14_10 = a[14]&b[10];
	assign in_15_10 = a[15]&b[10];
	assign in_16_10 = a[16]&b[10];
	assign in_17_10 = a[17]&b[10];
	assign in_18_10 = a[18]&b[10];
	assign in_19_10 = a[19]&b[10];
	assign in_20_10 = a[20]&b[10];
	assign in_21_10 = a[21]&b[10];
	assign in_22_10 = a[22]&b[10];
	assign in_23_10 = a[23]&b[10];
	assign in_24_10 = a[24]&b[10];
	assign in_25_10 = a[25]&b[10];
	assign in_26_10 = a[26]&b[10];
	assign in_27_10 = a[27]&b[10];
	assign in_28_10 = a[28]&b[10];
	assign in_29_10 = a[29]&b[10];
	assign in_30_10 = a[30]&b[10];
	assign in_31_10 = a[31]&b[10];
	assign in_0_11 = a[0]&b[11];
	assign in_1_11 = a[1]&b[11];
	assign in_2_11 = a[2]&b[11];
	assign in_3_11 = a[3]&b[11];
	assign in_4_11 = a[4]&b[11];
	assign in_5_11 = a[5]&b[11];
	assign in_6_11 = a[6]&b[11];
	assign in_7_11 = a[7]&b[11];
	assign in_8_11 = a[8]&b[11];
	assign in_9_11 = a[9]&b[11];
	assign in_10_11 = a[10]&b[11];
	assign in_11_11 = a[11]&b[11];
	assign in_12_11 = a[12]&b[11];
	assign in_13_11 = a[13]&b[11];
	assign in_14_11 = a[14]&b[11];
	assign in_15_11 = a[15]&b[11];
	assign in_16_11 = a[16]&b[11];
	assign in_17_11 = a[17]&b[11];
	assign in_18_11 = a[18]&b[11];
	assign in_19_11 = a[19]&b[11];
	assign in_20_11 = a[20]&b[11];
	assign in_21_11 = a[21]&b[11];
	assign in_22_11 = a[22]&b[11];
	assign in_23_11 = a[23]&b[11];
	assign in_24_11 = a[24]&b[11];
	assign in_25_11 = a[25]&b[11];
	assign in_26_11 = a[26]&b[11];
	assign in_27_11 = a[27]&b[11];
	assign in_28_11 = a[28]&b[11];
	assign in_29_11 = a[29]&b[11];
	assign in_30_11 = a[30]&b[11];
	assign in_31_11 = a[31]&b[11];
	assign in_0_12 = a[0]&b[12];
	assign in_1_12 = a[1]&b[12];
	assign in_2_12 = a[2]&b[12];
	assign in_3_12 = a[3]&b[12];
	assign in_4_12 = a[4]&b[12];
	assign in_5_12 = a[5]&b[12];
	assign in_6_12 = a[6]&b[12];
	assign in_7_12 = a[7]&b[12];
	assign in_8_12 = a[8]&b[12];
	assign in_9_12 = a[9]&b[12];
	assign in_10_12 = a[10]&b[12];
	assign in_11_12 = a[11]&b[12];
	assign in_12_12 = a[12]&b[12];
	assign in_13_12 = a[13]&b[12];
	assign in_14_12 = a[14]&b[12];
	assign in_15_12 = a[15]&b[12];
	assign in_16_12 = a[16]&b[12];
	assign in_17_12 = a[17]&b[12];
	assign in_18_12 = a[18]&b[12];
	assign in_19_12 = a[19]&b[12];
	assign in_20_12 = a[20]&b[12];
	assign in_21_12 = a[21]&b[12];
	assign in_22_12 = a[22]&b[12];
	assign in_23_12 = a[23]&b[12];
	assign in_24_12 = a[24]&b[12];
	assign in_25_12 = a[25]&b[12];
	assign in_26_12 = a[26]&b[12];
	assign in_27_12 = a[27]&b[12];
	assign in_28_12 = a[28]&b[12];
	assign in_29_12 = a[29]&b[12];
	assign in_30_12 = a[30]&b[12];
	assign in_31_12 = a[31]&b[12];
	assign in_0_13 = a[0]&b[13];
	assign in_1_13 = a[1]&b[13];
	assign in_2_13 = a[2]&b[13];
	assign in_3_13 = a[3]&b[13];
	assign in_4_13 = a[4]&b[13];
	assign in_5_13 = a[5]&b[13];
	assign in_6_13 = a[6]&b[13];
	assign in_7_13 = a[7]&b[13];
	assign in_8_13 = a[8]&b[13];
	assign in_9_13 = a[9]&b[13];
	assign in_10_13 = a[10]&b[13];
	assign in_11_13 = a[11]&b[13];
	assign in_12_13 = a[12]&b[13];
	assign in_13_13 = a[13]&b[13];
	assign in_14_13 = a[14]&b[13];
	assign in_15_13 = a[15]&b[13];
	assign in_16_13 = a[16]&b[13];
	assign in_17_13 = a[17]&b[13];
	assign in_18_13 = a[18]&b[13];
	assign in_19_13 = a[19]&b[13];
	assign in_20_13 = a[20]&b[13];
	assign in_21_13 = a[21]&b[13];
	assign in_22_13 = a[22]&b[13];
	assign in_23_13 = a[23]&b[13];
	assign in_24_13 = a[24]&b[13];
	assign in_25_13 = a[25]&b[13];
	assign in_26_13 = a[26]&b[13];
	assign in_27_13 = a[27]&b[13];
	assign in_28_13 = a[28]&b[13];
	assign in_29_13 = a[29]&b[13];
	assign in_30_13 = a[30]&b[13];
	assign in_31_13 = a[31]&b[13];
	assign in_0_14 = a[0]&b[14];
	assign in_1_14 = a[1]&b[14];
	assign in_2_14 = a[2]&b[14];
	assign in_3_14 = a[3]&b[14];
	assign in_4_14 = a[4]&b[14];
	assign in_5_14 = a[5]&b[14];
	assign in_6_14 = a[6]&b[14];
	assign in_7_14 = a[7]&b[14];
	assign in_8_14 = a[8]&b[14];
	assign in_9_14 = a[9]&b[14];
	assign in_10_14 = a[10]&b[14];
	assign in_11_14 = a[11]&b[14];
	assign in_12_14 = a[12]&b[14];
	assign in_13_14 = a[13]&b[14];
	assign in_14_14 = a[14]&b[14];
	assign in_15_14 = a[15]&b[14];
	assign in_16_14 = a[16]&b[14];
	assign in_17_14 = a[17]&b[14];
	assign in_18_14 = a[18]&b[14];
	assign in_19_14 = a[19]&b[14];
	assign in_20_14 = a[20]&b[14];
	assign in_21_14 = a[21]&b[14];
	assign in_22_14 = a[22]&b[14];
	assign in_23_14 = a[23]&b[14];
	assign in_24_14 = a[24]&b[14];
	assign in_25_14 = a[25]&b[14];
	assign in_26_14 = a[26]&b[14];
	assign in_27_14 = a[27]&b[14];
	assign in_28_14 = a[28]&b[14];
	assign in_29_14 = a[29]&b[14];
	assign in_30_14 = a[30]&b[14];
	assign in_31_14 = a[31]&b[14];
	assign in_0_15 = a[0]&b[15];
	assign in_1_15 = a[1]&b[15];
	assign in_2_15 = a[2]&b[15];
	assign in_3_15 = a[3]&b[15];
	assign in_4_15 = a[4]&b[15];
	assign in_5_15 = a[5]&b[15];
	assign in_6_15 = a[6]&b[15];
	assign in_7_15 = a[7]&b[15];
	assign in_8_15 = a[8]&b[15];
	assign in_9_15 = a[9]&b[15];
	assign in_10_15 = a[10]&b[15];
	assign in_11_15 = a[11]&b[15];
	assign in_12_15 = a[12]&b[15];
	assign in_13_15 = a[13]&b[15];
	assign in_14_15 = a[14]&b[15];
	assign in_15_15 = a[15]&b[15];
	assign in_16_15 = a[16]&b[15];
	assign in_17_15 = a[17]&b[15];
	assign in_18_15 = a[18]&b[15];
	assign in_19_15 = a[19]&b[15];
	assign in_20_15 = a[20]&b[15];
	assign in_21_15 = a[21]&b[15];
	assign in_22_15 = a[22]&b[15];
	assign in_23_15 = a[23]&b[15];
	assign in_24_15 = a[24]&b[15];
	assign in_25_15 = a[25]&b[15];
	assign in_26_15 = a[26]&b[15];
	assign in_27_15 = a[27]&b[15];
	assign in_28_15 = a[28]&b[15];
	assign in_29_15 = a[29]&b[15];
	assign in_30_15 = a[30]&b[15];
	assign in_31_15 = a[31]&b[15];
	assign in_0_16 = a[0]&b[16];
	assign in_1_16 = a[1]&b[16];
	assign in_2_16 = a[2]&b[16];
	assign in_3_16 = a[3]&b[16];
	assign in_4_16 = a[4]&b[16];
	assign in_5_16 = a[5]&b[16];
	assign in_6_16 = a[6]&b[16];
	assign in_7_16 = a[7]&b[16];
	assign in_8_16 = a[8]&b[16];
	assign in_9_16 = a[9]&b[16];
	assign in_10_16 = a[10]&b[16];
	assign in_11_16 = a[11]&b[16];
	assign in_12_16 = a[12]&b[16];
	assign in_13_16 = a[13]&b[16];
	assign in_14_16 = a[14]&b[16];
	assign in_15_16 = a[15]&b[16];
	assign in_16_16 = a[16]&b[16];
	assign in_17_16 = a[17]&b[16];
	assign in_18_16 = a[18]&b[16];
	assign in_19_16 = a[19]&b[16];
	assign in_20_16 = a[20]&b[16];
	assign in_21_16 = a[21]&b[16];
	assign in_22_16 = a[22]&b[16];
	assign in_23_16 = a[23]&b[16];
	assign in_24_16 = a[24]&b[16];
	assign in_25_16 = a[25]&b[16];
	assign in_26_16 = a[26]&b[16];
	assign in_27_16 = a[27]&b[16];
	assign in_28_16 = a[28]&b[16];
	assign in_29_16 = a[29]&b[16];
	assign in_30_16 = a[30]&b[16];
	assign in_31_16 = a[31]&b[16];
	assign in_0_17 = a[0]&b[17];
	assign in_1_17 = a[1]&b[17];
	assign in_2_17 = a[2]&b[17];
	assign in_3_17 = a[3]&b[17];
	assign in_4_17 = a[4]&b[17];
	assign in_5_17 = a[5]&b[17];
	assign in_6_17 = a[6]&b[17];
	assign in_7_17 = a[7]&b[17];
	assign in_8_17 = a[8]&b[17];
	assign in_9_17 = a[9]&b[17];
	assign in_10_17 = a[10]&b[17];
	assign in_11_17 = a[11]&b[17];
	assign in_12_17 = a[12]&b[17];
	assign in_13_17 = a[13]&b[17];
	assign in_14_17 = a[14]&b[17];
	assign in_15_17 = a[15]&b[17];
	assign in_16_17 = a[16]&b[17];
	assign in_17_17 = a[17]&b[17];
	assign in_18_17 = a[18]&b[17];
	assign in_19_17 = a[19]&b[17];
	assign in_20_17 = a[20]&b[17];
	assign in_21_17 = a[21]&b[17];
	assign in_22_17 = a[22]&b[17];
	assign in_23_17 = a[23]&b[17];
	assign in_24_17 = a[24]&b[17];
	assign in_25_17 = a[25]&b[17];
	assign in_26_17 = a[26]&b[17];
	assign in_27_17 = a[27]&b[17];
	assign in_28_17 = a[28]&b[17];
	assign in_29_17 = a[29]&b[17];
	assign in_30_17 = a[30]&b[17];
	assign in_31_17 = a[31]&b[17];
	assign in_0_18 = a[0]&b[18];
	assign in_1_18 = a[1]&b[18];
	assign in_2_18 = a[2]&b[18];
	assign in_3_18 = a[3]&b[18];
	assign in_4_18 = a[4]&b[18];
	assign in_5_18 = a[5]&b[18];
	assign in_6_18 = a[6]&b[18];
	assign in_7_18 = a[7]&b[18];
	assign in_8_18 = a[8]&b[18];
	assign in_9_18 = a[9]&b[18];
	assign in_10_18 = a[10]&b[18];
	assign in_11_18 = a[11]&b[18];
	assign in_12_18 = a[12]&b[18];
	assign in_13_18 = a[13]&b[18];
	assign in_14_18 = a[14]&b[18];
	assign in_15_18 = a[15]&b[18];
	assign in_16_18 = a[16]&b[18];
	assign in_17_18 = a[17]&b[18];
	assign in_18_18 = a[18]&b[18];
	assign in_19_18 = a[19]&b[18];
	assign in_20_18 = a[20]&b[18];
	assign in_21_18 = a[21]&b[18];
	assign in_22_18 = a[22]&b[18];
	assign in_23_18 = a[23]&b[18];
	assign in_24_18 = a[24]&b[18];
	assign in_25_18 = a[25]&b[18];
	assign in_26_18 = a[26]&b[18];
	assign in_27_18 = a[27]&b[18];
	assign in_28_18 = a[28]&b[18];
	assign in_29_18 = a[29]&b[18];
	assign in_30_18 = a[30]&b[18];
	assign in_31_18 = a[31]&b[18];
	assign in_0_19 = a[0]&b[19];
	assign in_1_19 = a[1]&b[19];
	assign in_2_19 = a[2]&b[19];
	assign in_3_19 = a[3]&b[19];
	assign in_4_19 = a[4]&b[19];
	assign in_5_19 = a[5]&b[19];
	assign in_6_19 = a[6]&b[19];
	assign in_7_19 = a[7]&b[19];
	assign in_8_19 = a[8]&b[19];
	assign in_9_19 = a[9]&b[19];
	assign in_10_19 = a[10]&b[19];
	assign in_11_19 = a[11]&b[19];
	assign in_12_19 = a[12]&b[19];
	assign in_13_19 = a[13]&b[19];
	assign in_14_19 = a[14]&b[19];
	assign in_15_19 = a[15]&b[19];
	assign in_16_19 = a[16]&b[19];
	assign in_17_19 = a[17]&b[19];
	assign in_18_19 = a[18]&b[19];
	assign in_19_19 = a[19]&b[19];
	assign in_20_19 = a[20]&b[19];
	assign in_21_19 = a[21]&b[19];
	assign in_22_19 = a[22]&b[19];
	assign in_23_19 = a[23]&b[19];
	assign in_24_19 = a[24]&b[19];
	assign in_25_19 = a[25]&b[19];
	assign in_26_19 = a[26]&b[19];
	assign in_27_19 = a[27]&b[19];
	assign in_28_19 = a[28]&b[19];
	assign in_29_19 = a[29]&b[19];
	assign in_30_19 = a[30]&b[19];
	assign in_31_19 = a[31]&b[19];
	assign in_0_20 = a[0]&b[20];
	assign in_1_20 = a[1]&b[20];
	assign in_2_20 = a[2]&b[20];
	assign in_3_20 = a[3]&b[20];
	assign in_4_20 = a[4]&b[20];
	assign in_5_20 = a[5]&b[20];
	assign in_6_20 = a[6]&b[20];
	assign in_7_20 = a[7]&b[20];
	assign in_8_20 = a[8]&b[20];
	assign in_9_20 = a[9]&b[20];
	assign in_10_20 = a[10]&b[20];
	assign in_11_20 = a[11]&b[20];
	assign in_12_20 = a[12]&b[20];
	assign in_13_20 = a[13]&b[20];
	assign in_14_20 = a[14]&b[20];
	assign in_15_20 = a[15]&b[20];
	assign in_16_20 = a[16]&b[20];
	assign in_17_20 = a[17]&b[20];
	assign in_18_20 = a[18]&b[20];
	assign in_19_20 = a[19]&b[20];
	assign in_20_20 = a[20]&b[20];
	assign in_21_20 = a[21]&b[20];
	assign in_22_20 = a[22]&b[20];
	assign in_23_20 = a[23]&b[20];
	assign in_24_20 = a[24]&b[20];
	assign in_25_20 = a[25]&b[20];
	assign in_26_20 = a[26]&b[20];
	assign in_27_20 = a[27]&b[20];
	assign in_28_20 = a[28]&b[20];
	assign in_29_20 = a[29]&b[20];
	assign in_30_20 = a[30]&b[20];
	assign in_31_20 = a[31]&b[20];
	assign in_0_21 = a[0]&b[21];
	assign in_1_21 = a[1]&b[21];
	assign in_2_21 = a[2]&b[21];
	assign in_3_21 = a[3]&b[21];
	assign in_4_21 = a[4]&b[21];
	assign in_5_21 = a[5]&b[21];
	assign in_6_21 = a[6]&b[21];
	assign in_7_21 = a[7]&b[21];
	assign in_8_21 = a[8]&b[21];
	assign in_9_21 = a[9]&b[21];
	assign in_10_21 = a[10]&b[21];
	assign in_11_21 = a[11]&b[21];
	assign in_12_21 = a[12]&b[21];
	assign in_13_21 = a[13]&b[21];
	assign in_14_21 = a[14]&b[21];
	assign in_15_21 = a[15]&b[21];
	assign in_16_21 = a[16]&b[21];
	assign in_17_21 = a[17]&b[21];
	assign in_18_21 = a[18]&b[21];
	assign in_19_21 = a[19]&b[21];
	assign in_20_21 = a[20]&b[21];
	assign in_21_21 = a[21]&b[21];
	assign in_22_21 = a[22]&b[21];
	assign in_23_21 = a[23]&b[21];
	assign in_24_21 = a[24]&b[21];
	assign in_25_21 = a[25]&b[21];
	assign in_26_21 = a[26]&b[21];
	assign in_27_21 = a[27]&b[21];
	assign in_28_21 = a[28]&b[21];
	assign in_29_21 = a[29]&b[21];
	assign in_30_21 = a[30]&b[21];
	assign in_31_21 = a[31]&b[21];
	assign in_0_22 = a[0]&b[22];
	assign in_1_22 = a[1]&b[22];
	assign in_2_22 = a[2]&b[22];
	assign in_3_22 = a[3]&b[22];
	assign in_4_22 = a[4]&b[22];
	assign in_5_22 = a[5]&b[22];
	assign in_6_22 = a[6]&b[22];
	assign in_7_22 = a[7]&b[22];
	assign in_8_22 = a[8]&b[22];
	assign in_9_22 = a[9]&b[22];
	assign in_10_22 = a[10]&b[22];
	assign in_11_22 = a[11]&b[22];
	assign in_12_22 = a[12]&b[22];
	assign in_13_22 = a[13]&b[22];
	assign in_14_22 = a[14]&b[22];
	assign in_15_22 = a[15]&b[22];
	assign in_16_22 = a[16]&b[22];
	assign in_17_22 = a[17]&b[22];
	assign in_18_22 = a[18]&b[22];
	assign in_19_22 = a[19]&b[22];
	assign in_20_22 = a[20]&b[22];
	assign in_21_22 = a[21]&b[22];
	assign in_22_22 = a[22]&b[22];
	assign in_23_22 = a[23]&b[22];
	assign in_24_22 = a[24]&b[22];
	assign in_25_22 = a[25]&b[22];
	assign in_26_22 = a[26]&b[22];
	assign in_27_22 = a[27]&b[22];
	assign in_28_22 = a[28]&b[22];
	assign in_29_22 = a[29]&b[22];
	assign in_30_22 = a[30]&b[22];
	assign in_31_22 = a[31]&b[22];
	assign in_0_23 = a[0]&b[23];
	assign in_1_23 = a[1]&b[23];
	assign in_2_23 = a[2]&b[23];
	assign in_3_23 = a[3]&b[23];
	assign in_4_23 = a[4]&b[23];
	assign in_5_23 = a[5]&b[23];
	assign in_6_23 = a[6]&b[23];
	assign in_7_23 = a[7]&b[23];
	assign in_8_23 = a[8]&b[23];
	assign in_9_23 = a[9]&b[23];
	assign in_10_23 = a[10]&b[23];
	assign in_11_23 = a[11]&b[23];
	assign in_12_23 = a[12]&b[23];
	assign in_13_23 = a[13]&b[23];
	assign in_14_23 = a[14]&b[23];
	assign in_15_23 = a[15]&b[23];
	assign in_16_23 = a[16]&b[23];
	assign in_17_23 = a[17]&b[23];
	assign in_18_23 = a[18]&b[23];
	assign in_19_23 = a[19]&b[23];
	assign in_20_23 = a[20]&b[23];
	assign in_21_23 = a[21]&b[23];
	assign in_22_23 = a[22]&b[23];
	assign in_23_23 = a[23]&b[23];
	assign in_24_23 = a[24]&b[23];
	assign in_25_23 = a[25]&b[23];
	assign in_26_23 = a[26]&b[23];
	assign in_27_23 = a[27]&b[23];
	assign in_28_23 = a[28]&b[23];
	assign in_29_23 = a[29]&b[23];
	assign in_30_23 = a[30]&b[23];
	assign in_31_23 = a[31]&b[23];
	assign in_0_24 = a[0]&b[24];
	assign in_1_24 = a[1]&b[24];
	assign in_2_24 = a[2]&b[24];
	assign in_3_24 = a[3]&b[24];
	assign in_4_24 = a[4]&b[24];
	assign in_5_24 = a[5]&b[24];
	assign in_6_24 = a[6]&b[24];
	assign in_7_24 = a[7]&b[24];
	assign in_8_24 = a[8]&b[24];
	assign in_9_24 = a[9]&b[24];
	assign in_10_24 = a[10]&b[24];
	assign in_11_24 = a[11]&b[24];
	assign in_12_24 = a[12]&b[24];
	assign in_13_24 = a[13]&b[24];
	assign in_14_24 = a[14]&b[24];
	assign in_15_24 = a[15]&b[24];
	assign in_16_24 = a[16]&b[24];
	assign in_17_24 = a[17]&b[24];
	assign in_18_24 = a[18]&b[24];
	assign in_19_24 = a[19]&b[24];
	assign in_20_24 = a[20]&b[24];
	assign in_21_24 = a[21]&b[24];
	assign in_22_24 = a[22]&b[24];
	assign in_23_24 = a[23]&b[24];
	assign in_24_24 = a[24]&b[24];
	assign in_25_24 = a[25]&b[24];
	assign in_26_24 = a[26]&b[24];
	assign in_27_24 = a[27]&b[24];
	assign in_28_24 = a[28]&b[24];
	assign in_29_24 = a[29]&b[24];
	assign in_30_24 = a[30]&b[24];
	assign in_31_24 = a[31]&b[24];
	assign in_0_25 = a[0]&b[25];
	assign in_1_25 = a[1]&b[25];
	assign in_2_25 = a[2]&b[25];
	assign in_3_25 = a[3]&b[25];
	assign in_4_25 = a[4]&b[25];
	assign in_5_25 = a[5]&b[25];
	assign in_6_25 = a[6]&b[25];
	assign in_7_25 = a[7]&b[25];
	assign in_8_25 = a[8]&b[25];
	assign in_9_25 = a[9]&b[25];
	assign in_10_25 = a[10]&b[25];
	assign in_11_25 = a[11]&b[25];
	assign in_12_25 = a[12]&b[25];
	assign in_13_25 = a[13]&b[25];
	assign in_14_25 = a[14]&b[25];
	assign in_15_25 = a[15]&b[25];
	assign in_16_25 = a[16]&b[25];
	assign in_17_25 = a[17]&b[25];
	assign in_18_25 = a[18]&b[25];
	assign in_19_25 = a[19]&b[25];
	assign in_20_25 = a[20]&b[25];
	assign in_21_25 = a[21]&b[25];
	assign in_22_25 = a[22]&b[25];
	assign in_23_25 = a[23]&b[25];
	assign in_24_25 = a[24]&b[25];
	assign in_25_25 = a[25]&b[25];
	assign in_26_25 = a[26]&b[25];
	assign in_27_25 = a[27]&b[25];
	assign in_28_25 = a[28]&b[25];
	assign in_29_25 = a[29]&b[25];
	assign in_30_25 = a[30]&b[25];
	assign in_31_25 = a[31]&b[25];
	assign in_0_26 = a[0]&b[26];
	assign in_1_26 = a[1]&b[26];
	assign in_2_26 = a[2]&b[26];
	assign in_3_26 = a[3]&b[26];
	assign in_4_26 = a[4]&b[26];
	assign in_5_26 = a[5]&b[26];
	assign in_6_26 = a[6]&b[26];
	assign in_7_26 = a[7]&b[26];
	assign in_8_26 = a[8]&b[26];
	assign in_9_26 = a[9]&b[26];
	assign in_10_26 = a[10]&b[26];
	assign in_11_26 = a[11]&b[26];
	assign in_12_26 = a[12]&b[26];
	assign in_13_26 = a[13]&b[26];
	assign in_14_26 = a[14]&b[26];
	assign in_15_26 = a[15]&b[26];
	assign in_16_26 = a[16]&b[26];
	assign in_17_26 = a[17]&b[26];
	assign in_18_26 = a[18]&b[26];
	assign in_19_26 = a[19]&b[26];
	assign in_20_26 = a[20]&b[26];
	assign in_21_26 = a[21]&b[26];
	assign in_22_26 = a[22]&b[26];
	assign in_23_26 = a[23]&b[26];
	assign in_24_26 = a[24]&b[26];
	assign in_25_26 = a[25]&b[26];
	assign in_26_26 = a[26]&b[26];
	assign in_27_26 = a[27]&b[26];
	assign in_28_26 = a[28]&b[26];
	assign in_29_26 = a[29]&b[26];
	assign in_30_26 = a[30]&b[26];
	assign in_31_26 = a[31]&b[26];
	assign in_0_27 = a[0]&b[27];
	assign in_1_27 = a[1]&b[27];
	assign in_2_27 = a[2]&b[27];
	assign in_3_27 = a[3]&b[27];
	assign in_4_27 = a[4]&b[27];
	assign in_5_27 = a[5]&b[27];
	assign in_6_27 = a[6]&b[27];
	assign in_7_27 = a[7]&b[27];
	assign in_8_27 = a[8]&b[27];
	assign in_9_27 = a[9]&b[27];
	assign in_10_27 = a[10]&b[27];
	assign in_11_27 = a[11]&b[27];
	assign in_12_27 = a[12]&b[27];
	assign in_13_27 = a[13]&b[27];
	assign in_14_27 = a[14]&b[27];
	assign in_15_27 = a[15]&b[27];
	assign in_16_27 = a[16]&b[27];
	assign in_17_27 = a[17]&b[27];
	assign in_18_27 = a[18]&b[27];
	assign in_19_27 = a[19]&b[27];
	assign in_20_27 = a[20]&b[27];
	assign in_21_27 = a[21]&b[27];
	assign in_22_27 = a[22]&b[27];
	assign in_23_27 = a[23]&b[27];
	assign in_24_27 = a[24]&b[27];
	assign in_25_27 = a[25]&b[27];
	assign in_26_27 = a[26]&b[27];
	assign in_27_27 = a[27]&b[27];
	assign in_28_27 = a[28]&b[27];
	assign in_29_27 = a[29]&b[27];
	assign in_30_27 = a[30]&b[27];
	assign in_31_27 = a[31]&b[27];
	assign in_0_28 = a[0]&b[28];
	assign in_1_28 = a[1]&b[28];
	assign in_2_28 = a[2]&b[28];
	assign in_3_28 = a[3]&b[28];
	assign in_4_28 = a[4]&b[28];
	assign in_5_28 = a[5]&b[28];
	assign in_6_28 = a[6]&b[28];
	assign in_7_28 = a[7]&b[28];
	assign in_8_28 = a[8]&b[28];
	assign in_9_28 = a[9]&b[28];
	assign in_10_28 = a[10]&b[28];
	assign in_11_28 = a[11]&b[28];
	assign in_12_28 = a[12]&b[28];
	assign in_13_28 = a[13]&b[28];
	assign in_14_28 = a[14]&b[28];
	assign in_15_28 = a[15]&b[28];
	assign in_16_28 = a[16]&b[28];
	assign in_17_28 = a[17]&b[28];
	assign in_18_28 = a[18]&b[28];
	assign in_19_28 = a[19]&b[28];
	assign in_20_28 = a[20]&b[28];
	assign in_21_28 = a[21]&b[28];
	assign in_22_28 = a[22]&b[28];
	assign in_23_28 = a[23]&b[28];
	assign in_24_28 = a[24]&b[28];
	assign in_25_28 = a[25]&b[28];
	assign in_26_28 = a[26]&b[28];
	assign in_27_28 = a[27]&b[28];
	assign in_28_28 = a[28]&b[28];
	assign in_29_28 = a[29]&b[28];
	assign in_30_28 = a[30]&b[28];
	assign in_31_28 = a[31]&b[28];
	assign in_0_29 = a[0]&b[29];
	assign in_1_29 = a[1]&b[29];
	assign in_2_29 = a[2]&b[29];
	assign in_3_29 = a[3]&b[29];
	assign in_4_29 = a[4]&b[29];
	assign in_5_29 = a[5]&b[29];
	assign in_6_29 = a[6]&b[29];
	assign in_7_29 = a[7]&b[29];
	assign in_8_29 = a[8]&b[29];
	assign in_9_29 = a[9]&b[29];
	assign in_10_29 = a[10]&b[29];
	assign in_11_29 = a[11]&b[29];
	assign in_12_29 = a[12]&b[29];
	assign in_13_29 = a[13]&b[29];
	assign in_14_29 = a[14]&b[29];
	assign in_15_29 = a[15]&b[29];
	assign in_16_29 = a[16]&b[29];
	assign in_17_29 = a[17]&b[29];
	assign in_18_29 = a[18]&b[29];
	assign in_19_29 = a[19]&b[29];
	assign in_20_29 = a[20]&b[29];
	assign in_21_29 = a[21]&b[29];
	assign in_22_29 = a[22]&b[29];
	assign in_23_29 = a[23]&b[29];
	assign in_24_29 = a[24]&b[29];
	assign in_25_29 = a[25]&b[29];
	assign in_26_29 = a[26]&b[29];
	assign in_27_29 = a[27]&b[29];
	assign in_28_29 = a[28]&b[29];
	assign in_29_29 = a[29]&b[29];
	assign in_30_29 = a[30]&b[29];
	assign in_31_29 = a[31]&b[29];
	assign in_0_30 = a[0]&b[30];
	assign in_1_30 = a[1]&b[30];
	assign in_2_30 = a[2]&b[30];
	assign in_3_30 = a[3]&b[30];
	assign in_4_30 = a[4]&b[30];
	assign in_5_30 = a[5]&b[30];
	assign in_6_30 = a[6]&b[30];
	assign in_7_30 = a[7]&b[30];
	assign in_8_30 = a[8]&b[30];
	assign in_9_30 = a[9]&b[30];
	assign in_10_30 = a[10]&b[30];
	assign in_11_30 = a[11]&b[30];
	assign in_12_30 = a[12]&b[30];
	assign in_13_30 = a[13]&b[30];
	assign in_14_30 = a[14]&b[30];
	assign in_15_30 = a[15]&b[30];
	assign in_16_30 = a[16]&b[30];
	assign in_17_30 = a[17]&b[30];
	assign in_18_30 = a[18]&b[30];
	assign in_19_30 = a[19]&b[30];
	assign in_20_30 = a[20]&b[30];
	assign in_21_30 = a[21]&b[30];
	assign in_22_30 = a[22]&b[30];
	assign in_23_30 = a[23]&b[30];
	assign in_24_30 = a[24]&b[30];
	assign in_25_30 = a[25]&b[30];
	assign in_26_30 = a[26]&b[30];
	assign in_27_30 = a[27]&b[30];
	assign in_28_30 = a[28]&b[30];
	assign in_29_30 = a[29]&b[30];
	assign in_30_30 = a[30]&b[30];
	assign in_31_30 = a[31]&b[30];
	assign in_0_31 = a[0]&b[31];
	assign in_1_31 = a[1]&b[31];
	assign in_2_31 = a[2]&b[31];
	assign in_3_31 = a[3]&b[31];
	assign in_4_31 = a[4]&b[31];
	assign in_5_31 = a[5]&b[31];
	assign in_6_31 = a[6]&b[31];
	assign in_7_31 = a[7]&b[31];
	assign in_8_31 = a[8]&b[31];
	assign in_9_31 = a[9]&b[31];
	assign in_10_31 = a[10]&b[31];
	assign in_11_31 = a[11]&b[31];
	assign in_12_31 = a[12]&b[31];
	assign in_13_31 = a[13]&b[31];
	assign in_14_31 = a[14]&b[31];
	assign in_15_31 = a[15]&b[31];
	assign in_16_31 = a[16]&b[31];
	assign in_17_31 = a[17]&b[31];
	assign in_18_31 = a[18]&b[31];
	assign in_19_31 = a[19]&b[31];
	assign in_20_31 = a[20]&b[31];
	assign in_21_31 = a[21]&b[31];
	assign in_22_31 = a[22]&b[31];
	assign in_23_31 = a[23]&b[31];
	assign in_24_31 = a[24]&b[31];
	assign in_25_31 = a[25]&b[31];
	assign in_26_31 = a[26]&b[31];
	assign in_27_31 = a[27]&b[31];
	assign in_28_31 = a[28]&b[31];
	assign in_29_31 = a[29]&b[31];
	assign in_30_31 = a[30]&b[31];
	assign in_31_31 = a[31]&b[31];

	logic fs0, fc0;
	FA fa0 (.a(in_0_2), .b(in_1_1), .c_in(in_2_0), .s(fs0), .c_out(fc0));

	logic hs3, hc3;
	HA ha3 (.a(in_0_3), .b(in_1_2), .s(hs3), .c_out(hc3));

	logic fs1, fc1;
	FA fa1 (.a(in_2_1), .b(in_3_0), .c_in(hs3), .s(fs1), .c_out(fc1));

	logic hs4, hc4;
	HA ha4 (.a(in_0_4), .b(in_1_3), .s(hs4), .c_out(hc4));

	logic fs2, fc2;
	FA fa2 (.a(in_2_2), .b(in_3_1), .c_in(in_4_0), .s(fs2), .c_out(fc2));

	logic fs3, fc3;
	FA fa3 (.a(hc3), .b(hs4), .c_in(fs2), .s(fs3), .c_out(fc3));

	logic hs5, hc5;
	HA ha5 (.a(in_0_5), .b(in_1_4), .s(hs5), .c_out(hc5));

	logic fs4, fc4;
	FA fa4 (.a(in_2_3), .b(in_3_2), .c_in(in_4_1), .s(fs4), .c_out(fc4));

	logic fs5, fc5;
	FA fa5 (.a(in_5_0), .b(hc4), .c_in(hs5), .s(fs5), .c_out(fc5));

	logic fs6, fc6;
	FA fa6 (.a(fc2), .b(fs4), .c_in(fs5), .s(fs6), .c_out(fc6));

	logic hs6, hc6;
	HA ha6 (.a(in_0_6), .b(in_1_5), .s(hs6), .c_out(hc6));

	logic fs7, fc7;
	FA fa7 (.a(in_2_4), .b(in_3_3), .c_in(in_4_2), .s(fs7), .c_out(fc7));

	logic fs8, fc8;
	FA fa8 (.a(in_5_1), .b(in_6_0), .c_in(hc5), .s(fs8), .c_out(fc8));

	logic fs9, fc9;
	FA fa9 (.a(hs6), .b(fc4), .c_in(fc5), .s(fs9), .c_out(fc9));

	logic fs10, fc10;
	FA fa10 (.a(fs7), .b(fs8), .c_in(fs9), .s(fs10), .c_out(fc10));

	logic hs7, hc7;
	HA ha7 (.a(in_0_7), .b(in_1_6), .s(hs7), .c_out(hc7));

	logic fs11, fc11;
	FA fa11 (.a(in_2_5), .b(in_3_4), .c_in(in_4_3), .s(fs11), .c_out(fc11));

	logic fs12, fc12;
	FA fa12 (.a(in_5_2), .b(in_6_1), .c_in(in_7_0), .s(fs12), .c_out(fc12));

	logic fs13, fc13;
	FA fa13 (.a(hc6), .b(hs7), .c_in(fc7), .s(fs13), .c_out(fc13));

	logic fs14, fc14;
	FA fa14 (.a(fc8), .b(fs11), .c_in(fs12), .s(fs14), .c_out(fc14));

	logic fs15, fc15;
	FA fa15 (.a(fc9), .b(fs13), .c_in(fs14), .s(fs15), .c_out(fc15));

	logic hs8, hc8;
	HA ha8 (.a(in_0_8), .b(in_1_7), .s(hs8), .c_out(hc8));

	logic fs16, fc16;
	FA fa16 (.a(in_2_6), .b(in_3_5), .c_in(in_4_4), .s(fs16), .c_out(fc16));

	logic fs17, fc17;
	FA fa17 (.a(in_5_3), .b(in_6_2), .c_in(in_7_1), .s(fs17), .c_out(fc17));

	logic fs18, fc18;
	FA fa18 (.a(in_8_0), .b(hc7), .c_in(hs8), .s(fs18), .c_out(fc18));

	logic fs19, fc19;
	FA fa19 (.a(fc11), .b(fc12), .c_in(fc13), .s(fs19), .c_out(fc19));

	logic fs20, fc20;
	FA fa20 (.a(fs16), .b(fs17), .c_in(fs18), .s(fs20), .c_out(fc20));

	logic fs21, fc21;
	FA fa21 (.a(fc14), .b(fs19), .c_in(fs20), .s(fs21), .c_out(fc21));

	logic hs9, hc9;
	HA ha9 (.a(in_0_9), .b(in_1_8), .s(hs9), .c_out(hc9));

	logic fs22, fc22;
	FA fa22 (.a(in_2_7), .b(in_3_6), .c_in(in_4_5), .s(fs22), .c_out(fc22));

	logic fs23, fc23;
	FA fa23 (.a(in_5_4), .b(in_6_3), .c_in(in_7_2), .s(fs23), .c_out(fc23));

	logic fs24, fc24;
	FA fa24 (.a(in_8_1), .b(in_9_0), .c_in(hc8), .s(fs24), .c_out(fc24));

	logic fs25, fc25;
	FA fa25 (.a(hs9), .b(fc16), .c_in(fc17), .s(fs25), .c_out(fc25));

	logic fs26, fc26;
	FA fa26 (.a(fc18), .b(fs22), .c_in(fs23), .s(fs26), .c_out(fc26));

	logic fs27, fc27;
	FA fa27 (.a(fs24), .b(fc19), .c_in(fc20), .s(fs27), .c_out(fc27));

	logic fs28, fc28;
	FA fa28 (.a(fs25), .b(fs26), .c_in(fs27), .s(fs28), .c_out(fc28));

	logic hs10, hc10;
	HA ha10 (.a(in_0_10), .b(in_1_9), .s(hs10), .c_out(hc10));

	logic fs29, fc29;
	FA fa29 (.a(in_2_8), .b(in_3_7), .c_in(in_4_6), .s(fs29), .c_out(fc29));

	logic fs30, fc30;
	FA fa30 (.a(in_5_5), .b(in_6_4), .c_in(in_7_3), .s(fs30), .c_out(fc30));

	logic fs31, fc31;
	FA fa31 (.a(in_8_2), .b(in_9_1), .c_in(in_10_0), .s(fs31), .c_out(fc31));

	logic fs32, fc32;
	FA fa32 (.a(hc9), .b(hs10), .c_in(fc22), .s(fs32), .c_out(fc32));

	logic fs33, fc33;
	FA fa33 (.a(fc23), .b(fc24), .c_in(fs29), .s(fs33), .c_out(fc33));

	logic fs34, fc34;
	FA fa34 (.a(fs30), .b(fs31), .c_in(fc25), .s(fs34), .c_out(fc34));

	logic fs35, fc35;
	FA fa35 (.a(fs32), .b(fc26), .c_in(fs33), .s(fs35), .c_out(fc35));

	logic fs36, fc36;
	FA fa36 (.a(fc27), .b(fs34), .c_in(fs35), .s(fs36), .c_out(fc36));

	logic hs11, hc11;
	HA ha11 (.a(in_0_11), .b(in_1_10), .s(hs11), .c_out(hc11));

	logic fs37, fc37;
	FA fa37 (.a(in_2_9), .b(in_3_8), .c_in(in_4_7), .s(fs37), .c_out(fc37));

	logic fs38, fc38;
	FA fa38 (.a(in_5_6), .b(in_6_5), .c_in(in_7_4), .s(fs38), .c_out(fc38));

	logic fs39, fc39;
	FA fa39 (.a(in_8_3), .b(in_9_2), .c_in(in_10_1), .s(fs39), .c_out(fc39));

	logic fs40, fc40;
	FA fa40 (.a(in_11_0), .b(hc10), .c_in(hs11), .s(fs40), .c_out(fc40));

	logic fs41, fc41;
	FA fa41 (.a(fc29), .b(fc30), .c_in(fc31), .s(fs41), .c_out(fc41));

	logic fs42, fc42;
	FA fa42 (.a(fc32), .b(fs37), .c_in(fs38), .s(fs42), .c_out(fc42));

	logic fs43, fc43;
	FA fa43 (.a(fs39), .b(fs40), .c_in(fc33), .s(fs43), .c_out(fc43));

	logic fs44, fc44;
	FA fa44 (.a(fc34), .b(fs41), .c_in(fs42), .s(fs44), .c_out(fc44));

	logic fs45, fc45;
	FA fa45 (.a(fs43), .b(fc35), .c_in(fs44), .s(fs45), .c_out(fc45));

	logic hs12, hc12;
	HA ha12 (.a(in_0_12), .b(in_1_11), .s(hs12), .c_out(hc12));

	logic fs46, fc46;
	FA fa46 (.a(in_2_10), .b(in_3_9), .c_in(in_4_8), .s(fs46), .c_out(fc46));

	logic fs47, fc47;
	FA fa47 (.a(in_5_7), .b(in_6_6), .c_in(in_7_5), .s(fs47), .c_out(fc47));

	logic fs48, fc48;
	FA fa48 (.a(in_8_4), .b(in_9_3), .c_in(in_10_2), .s(fs48), .c_out(fc48));

	logic fs49, fc49;
	FA fa49 (.a(in_11_1), .b(in_12_0), .c_in(hc11), .s(fs49), .c_out(fc49));

	logic fs50, fc50;
	FA fa50 (.a(hs12), .b(fc37), .c_in(fc38), .s(fs50), .c_out(fc50));

	logic fs51, fc51;
	FA fa51 (.a(fc39), .b(fc40), .c_in(fs46), .s(fs51), .c_out(fc51));

	logic fs52, fc52;
	FA fa52 (.a(fs47), .b(fs48), .c_in(fs49), .s(fs52), .c_out(fc52));

	logic fs53, fc53;
	FA fa53 (.a(fc41), .b(fc42), .c_in(fs50), .s(fs53), .c_out(fc53));

	logic fs54, fc54;
	FA fa54 (.a(fc43), .b(fs51), .c_in(fs52), .s(fs54), .c_out(fc54));

	logic fs55, fc55;
	FA fa55 (.a(fc44), .b(fs53), .c_in(fs54), .s(fs55), .c_out(fc55));

	logic hs13, hc13;
	HA ha13 (.a(in_0_13), .b(in_1_12), .s(hs13), .c_out(hc13));

	logic fs56, fc56;
	FA fa56 (.a(in_2_11), .b(in_3_10), .c_in(in_4_9), .s(fs56), .c_out(fc56));

	logic fs57, fc57;
	FA fa57 (.a(in_5_8), .b(in_6_7), .c_in(in_7_6), .s(fs57), .c_out(fc57));

	logic fs58, fc58;
	FA fa58 (.a(in_8_5), .b(in_9_4), .c_in(in_10_3), .s(fs58), .c_out(fc58));

	logic fs59, fc59;
	FA fa59 (.a(in_11_2), .b(in_12_1), .c_in(in_13_0), .s(fs59), .c_out(fc59));

	logic fs60, fc60;
	FA fa60 (.a(hc12), .b(hs13), .c_in(fc46), .s(fs60), .c_out(fc60));

	logic fs61, fc61;
	FA fa61 (.a(fc47), .b(fc48), .c_in(fc49), .s(fs61), .c_out(fc61));

	logic fs62, fc62;
	FA fa62 (.a(fs56), .b(fs57), .c_in(fs58), .s(fs62), .c_out(fc62));

	logic fs63, fc63;
	FA fa63 (.a(fs59), .b(fc50), .c_in(fs60), .s(fs63), .c_out(fc63));

	logic fs64, fc64;
	FA fa64 (.a(fc51), .b(fc52), .c_in(fs61), .s(fs64), .c_out(fc64));

	logic fs65, fc65;
	FA fa65 (.a(fs62), .b(fc53), .c_in(fs63), .s(fs65), .c_out(fc65));

	logic fs66, fc66;
	FA fa66 (.a(fc54), .b(fs64), .c_in(fs65), .s(fs66), .c_out(fc66));

	logic hs14, hc14;
	HA ha14 (.a(in_0_14), .b(in_1_13), .s(hs14), .c_out(hc14));

	logic fs67, fc67;
	FA fa67 (.a(in_2_12), .b(in_3_11), .c_in(in_4_10), .s(fs67), .c_out(fc67));

	logic fs68, fc68;
	FA fa68 (.a(in_5_9), .b(in_6_8), .c_in(in_7_7), .s(fs68), .c_out(fc68));

	logic fs69, fc69;
	FA fa69 (.a(in_8_6), .b(in_9_5), .c_in(in_10_4), .s(fs69), .c_out(fc69));

	logic fs70, fc70;
	FA fa70 (.a(in_11_3), .b(in_12_2), .c_in(in_13_1), .s(fs70), .c_out(fc70));

	logic fs71, fc71;
	FA fa71 (.a(in_14_0), .b(hc13), .c_in(hs14), .s(fs71), .c_out(fc71));

	logic fs72, fc72;
	FA fa72 (.a(fc56), .b(fc57), .c_in(fc58), .s(fs72), .c_out(fc72));

	logic fs73, fc73;
	FA fa73 (.a(fc59), .b(fc60), .c_in(fs67), .s(fs73), .c_out(fc73));

	logic fs74, fc74;
	FA fa74 (.a(fs68), .b(fs69), .c_in(fs70), .s(fs74), .c_out(fc74));

	logic fs75, fc75;
	FA fa75 (.a(fs71), .b(fc61), .c_in(fc62), .s(fs75), .c_out(fc75));

	logic fs76, fc76;
	FA fa76 (.a(fs72), .b(fc63), .c_in(fs73), .s(fs76), .c_out(fc76));

	logic fs77, fc77;
	FA fa77 (.a(fs74), .b(fc64), .c_in(fs75), .s(fs77), .c_out(fc77));

	logic fs78, fc78;
	FA fa78 (.a(fc65), .b(fs76), .c_in(fs77), .s(fs78), .c_out(fc78));

	logic hs15, hc15;
	HA ha15 (.a(in_0_15), .b(in_1_14), .s(hs15), .c_out(hc15));

	logic fs79, fc79;
	FA fa79 (.a(in_2_13), .b(in_3_12), .c_in(in_4_11), .s(fs79), .c_out(fc79));

	logic fs80, fc80;
	FA fa80 (.a(in_5_10), .b(in_6_9), .c_in(in_7_8), .s(fs80), .c_out(fc80));

	logic fs81, fc81;
	FA fa81 (.a(in_8_7), .b(in_9_6), .c_in(in_10_5), .s(fs81), .c_out(fc81));

	logic fs82, fc82;
	FA fa82 (.a(in_11_4), .b(in_12_3), .c_in(in_13_2), .s(fs82), .c_out(fc82));

	logic fs83, fc83;
	FA fa83 (.a(in_14_1), .b(in_15_0), .c_in(hc14), .s(fs83), .c_out(fc83));

	logic fs84, fc84;
	FA fa84 (.a(hs15), .b(fc67), .c_in(fc68), .s(fs84), .c_out(fc84));

	logic fs85, fc85;
	FA fa85 (.a(fc69), .b(fc70), .c_in(fc71), .s(fs85), .c_out(fc85));

	logic fs86, fc86;
	FA fa86 (.a(fs79), .b(fs80), .c_in(fs81), .s(fs86), .c_out(fc86));

	logic fs87, fc87;
	FA fa87 (.a(fs82), .b(fs83), .c_in(fc72), .s(fs87), .c_out(fc87));

	logic fs88, fc88;
	FA fa88 (.a(fc73), .b(fc74), .c_in(fs84), .s(fs88), .c_out(fc88));

	logic fs89, fc89;
	FA fa89 (.a(fs85), .b(fc75), .c_in(fs86), .s(fs89), .c_out(fc89));

	logic fs90, fc90;
	FA fa90 (.a(fs87), .b(fc76), .c_in(fs88), .s(fs90), .c_out(fc90));

	logic fs91, fc91;
	FA fa91 (.a(fc77), .b(fs89), .c_in(fs90), .s(fs91), .c_out(fc91));

	logic hs16, hc16;
	HA ha16 (.a(in_0_16), .b(in_1_15), .s(hs16), .c_out(hc16));

	logic fs92, fc92;
	FA fa92 (.a(in_2_14), .b(in_3_13), .c_in(in_4_12), .s(fs92), .c_out(fc92));

	logic fs93, fc93;
	FA fa93 (.a(in_5_11), .b(in_6_10), .c_in(in_7_9), .s(fs93), .c_out(fc93));

	logic fs94, fc94;
	FA fa94 (.a(in_8_8), .b(in_9_7), .c_in(in_10_6), .s(fs94), .c_out(fc94));

	logic fs95, fc95;
	FA fa95 (.a(in_11_5), .b(in_12_4), .c_in(in_13_3), .s(fs95), .c_out(fc95));

	logic fs96, fc96;
	FA fa96 (.a(in_14_2), .b(in_15_1), .c_in(in_16_0), .s(fs96), .c_out(fc96));

	logic fs97, fc97;
	FA fa97 (.a(hc15), .b(hs16), .c_in(fc79), .s(fs97), .c_out(fc97));

	logic fs98, fc98;
	FA fa98 (.a(fc80), .b(fc81), .c_in(fc82), .s(fs98), .c_out(fc98));

	logic fs99, fc99;
	FA fa99 (.a(fc83), .b(fs92), .c_in(fs93), .s(fs99), .c_out(fc99));

	logic fs100, fc100;
	FA fa100 (.a(fs94), .b(fs95), .c_in(fs96), .s(fs100), .c_out(fc100));

	logic fs101, fc101;
	FA fa101 (.a(fc84), .b(fc85), .c_in(fs97), .s(fs101), .c_out(fc101));

	logic fs102, fc102;
	FA fa102 (.a(fc86), .b(fc87), .c_in(fs98), .s(fs102), .c_out(fc102));

	logic fs103, fc103;
	FA fa103 (.a(fs99), .b(fs100), .c_in(fc88), .s(fs103), .c_out(fc103));

	logic fs104, fc104;
	FA fa104 (.a(fs101), .b(fc89), .c_in(fs102), .s(fs104), .c_out(fc104));

	logic fs105, fc105;
	FA fa105 (.a(fs103), .b(fc90), .c_in(fs104), .s(fs105), .c_out(fc105));

	logic hs17, hc17;
	HA ha17 (.a(in_0_17), .b(in_1_16), .s(hs17), .c_out(hc17));

	logic fs106, fc106;
	FA fa106 (.a(in_2_15), .b(in_3_14), .c_in(in_4_13), .s(fs106), .c_out(fc106));

	logic fs107, fc107;
	FA fa107 (.a(in_5_12), .b(in_6_11), .c_in(in_7_10), .s(fs107), .c_out(fc107));

	logic fs108, fc108;
	FA fa108 (.a(in_8_9), .b(in_9_8), .c_in(in_10_7), .s(fs108), .c_out(fc108));

	logic fs109, fc109;
	FA fa109 (.a(in_11_6), .b(in_12_5), .c_in(in_13_4), .s(fs109), .c_out(fc109));

	logic fs110, fc110;
	FA fa110 (.a(in_14_3), .b(in_15_2), .c_in(in_16_1), .s(fs110), .c_out(fc110));

	logic fs111, fc111;
	FA fa111 (.a(in_17_0), .b(hc16), .c_in(hs17), .s(fs111), .c_out(fc111));

	logic fs112, fc112;
	FA fa112 (.a(fc92), .b(fc93), .c_in(fc94), .s(fs112), .c_out(fc112));

	logic fs113, fc113;
	FA fa113 (.a(fc95), .b(fc96), .c_in(fc97), .s(fs113), .c_out(fc113));

	logic fs114, fc114;
	FA fa114 (.a(fs106), .b(fs107), .c_in(fs108), .s(fs114), .c_out(fc114));

	logic fs115, fc115;
	FA fa115 (.a(fs109), .b(fs110), .c_in(fs111), .s(fs115), .c_out(fc115));

	logic fs116, fc116;
	FA fa116 (.a(fc98), .b(fc99), .c_in(fc100), .s(fs116), .c_out(fc116));

	logic fs117, fc117;
	FA fa117 (.a(fs112), .b(fs113), .c_in(fc101), .s(fs117), .c_out(fc117));

	logic fs118, fc118;
	FA fa118 (.a(fs114), .b(fs115), .c_in(fc102), .s(fs118), .c_out(fc118));

	logic fs119, fc119;
	FA fa119 (.a(fc103), .b(fs116), .c_in(fs117), .s(fs119), .c_out(fc119));

	logic fs120, fc120;
	FA fa120 (.a(fs118), .b(fc104), .c_in(fs119), .s(fs120), .c_out(fc120));

	logic hs18, hc18;
	HA ha18 (.a(in_0_18), .b(in_1_17), .s(hs18), .c_out(hc18));

	logic fs121, fc121;
	FA fa121 (.a(in_2_16), .b(in_3_15), .c_in(in_4_14), .s(fs121), .c_out(fc121));

	logic fs122, fc122;
	FA fa122 (.a(in_5_13), .b(in_6_12), .c_in(in_7_11), .s(fs122), .c_out(fc122));

	logic fs123, fc123;
	FA fa123 (.a(in_8_10), .b(in_9_9), .c_in(in_10_8), .s(fs123), .c_out(fc123));

	logic fs124, fc124;
	FA fa124 (.a(in_11_7), .b(in_12_6), .c_in(in_13_5), .s(fs124), .c_out(fc124));

	logic fs125, fc125;
	FA fa125 (.a(in_14_4), .b(in_15_3), .c_in(in_16_2), .s(fs125), .c_out(fc125));

	logic fs126, fc126;
	FA fa126 (.a(in_17_1), .b(in_18_0), .c_in(hc17), .s(fs126), .c_out(fc126));

	logic fs127, fc127;
	FA fa127 (.a(hs18), .b(fc106), .c_in(fc107), .s(fs127), .c_out(fc127));

	logic fs128, fc128;
	FA fa128 (.a(fc108), .b(fc109), .c_in(fc110), .s(fs128), .c_out(fc128));

	logic fs129, fc129;
	FA fa129 (.a(fc111), .b(fs121), .c_in(fs122), .s(fs129), .c_out(fc129));

	logic fs130, fc130;
	FA fa130 (.a(fs123), .b(fs124), .c_in(fs125), .s(fs130), .c_out(fc130));

	logic fs131, fc131;
	FA fa131 (.a(fs126), .b(fc112), .c_in(fc113), .s(fs131), .c_out(fc131));

	logic fs132, fc132;
	FA fa132 (.a(fc114), .b(fc115), .c_in(fs127), .s(fs132), .c_out(fc132));

	logic fs133, fc133;
	FA fa133 (.a(fs128), .b(fs129), .c_in(fs130), .s(fs133), .c_out(fc133));

	logic fs134, fc134;
	FA fa134 (.a(fc116), .b(fc117), .c_in(fs131), .s(fs134), .c_out(fc134));

	logic fs135, fc135;
	FA fa135 (.a(fc118), .b(fs132), .c_in(fs133), .s(fs135), .c_out(fc135));

	logic fs136, fc136;
	FA fa136 (.a(fc119), .b(fs134), .c_in(fs135), .s(fs136), .c_out(fc136));

	logic hs19, hc19;
	HA ha19 (.a(in_0_19), .b(in_1_18), .s(hs19), .c_out(hc19));

	logic fs137, fc137;
	FA fa137 (.a(in_2_17), .b(in_3_16), .c_in(in_4_15), .s(fs137), .c_out(fc137));

	logic fs138, fc138;
	FA fa138 (.a(in_5_14), .b(in_6_13), .c_in(in_7_12), .s(fs138), .c_out(fc138));

	logic fs139, fc139;
	FA fa139 (.a(in_8_11), .b(in_9_10), .c_in(in_10_9), .s(fs139), .c_out(fc139));

	logic fs140, fc140;
	FA fa140 (.a(in_11_8), .b(in_12_7), .c_in(in_13_6), .s(fs140), .c_out(fc140));

	logic fs141, fc141;
	FA fa141 (.a(in_14_5), .b(in_15_4), .c_in(in_16_3), .s(fs141), .c_out(fc141));

	logic fs142, fc142;
	FA fa142 (.a(in_17_2), .b(in_18_1), .c_in(in_19_0), .s(fs142), .c_out(fc142));

	logic fs143, fc143;
	FA fa143 (.a(hc18), .b(hs19), .c_in(fc121), .s(fs143), .c_out(fc143));

	logic fs144, fc144;
	FA fa144 (.a(fc122), .b(fc123), .c_in(fc124), .s(fs144), .c_out(fc144));

	logic fs145, fc145;
	FA fa145 (.a(fc125), .b(fc126), .c_in(fs137), .s(fs145), .c_out(fc145));

	logic fs146, fc146;
	FA fa146 (.a(fs138), .b(fs139), .c_in(fs140), .s(fs146), .c_out(fc146));

	logic fs147, fc147;
	FA fa147 (.a(fs141), .b(fs142), .c_in(fc127), .s(fs147), .c_out(fc147));

	logic fs148, fc148;
	FA fa148 (.a(fc128), .b(fs143), .c_in(fc129), .s(fs148), .c_out(fc148));

	logic fs149, fc149;
	FA fa149 (.a(fc130), .b(fs144), .c_in(fs145), .s(fs149), .c_out(fc149));

	logic fs150, fc150;
	FA fa150 (.a(fc131), .b(fs146), .c_in(fs147), .s(fs150), .c_out(fc150));

	logic fs151, fc151;
	FA fa151 (.a(fc132), .b(fs148), .c_in(fc133), .s(fs151), .c_out(fc151));

	logic fs152, fc152;
	FA fa152 (.a(fs149), .b(fc134), .c_in(fs150), .s(fs152), .c_out(fc152));

	logic fs153, fc153;
	FA fa153 (.a(fc135), .b(fs151), .c_in(fs152), .s(fs153), .c_out(fc153));

	logic hs20, hc20;
	HA ha20 (.a(in_0_20), .b(in_1_19), .s(hs20), .c_out(hc20));

	logic fs154, fc154;
	FA fa154 (.a(in_2_18), .b(in_3_17), .c_in(in_4_16), .s(fs154), .c_out(fc154));

	logic fs155, fc155;
	FA fa155 (.a(in_5_15), .b(in_6_14), .c_in(in_7_13), .s(fs155), .c_out(fc155));

	logic fs156, fc156;
	FA fa156 (.a(in_8_12), .b(in_9_11), .c_in(in_10_10), .s(fs156), .c_out(fc156));

	logic fs157, fc157;
	FA fa157 (.a(in_11_9), .b(in_12_8), .c_in(in_13_7), .s(fs157), .c_out(fc157));

	logic fs158, fc158;
	FA fa158 (.a(in_14_6), .b(in_15_5), .c_in(in_16_4), .s(fs158), .c_out(fc158));

	logic fs159, fc159;
	FA fa159 (.a(in_17_3), .b(in_18_2), .c_in(in_19_1), .s(fs159), .c_out(fc159));

	logic fs160, fc160;
	FA fa160 (.a(in_20_0), .b(hc19), .c_in(hs20), .s(fs160), .c_out(fc160));

	logic fs161, fc161;
	FA fa161 (.a(fc137), .b(fc138), .c_in(fc139), .s(fs161), .c_out(fc161));

	logic fs162, fc162;
	FA fa162 (.a(fc140), .b(fc141), .c_in(fc142), .s(fs162), .c_out(fc162));

	logic fs163, fc163;
	FA fa163 (.a(fc143), .b(fs154), .c_in(fs155), .s(fs163), .c_out(fc163));

	logic fs164, fc164;
	FA fa164 (.a(fs156), .b(fs157), .c_in(fs158), .s(fs164), .c_out(fc164));

	logic fs165, fc165;
	FA fa165 (.a(fs159), .b(fs160), .c_in(fc144), .s(fs165), .c_out(fc165));

	logic fs166, fc166;
	FA fa166 (.a(fc145), .b(fc146), .c_in(fc147), .s(fs166), .c_out(fc166));

	logic fs167, fc167;
	FA fa167 (.a(fs161), .b(fs162), .c_in(fc148), .s(fs167), .c_out(fc167));

	logic fs168, fc168;
	FA fa168 (.a(fs163), .b(fs164), .c_in(fs165), .s(fs168), .c_out(fc168));

	logic fs169, fc169;
	FA fa169 (.a(fc149), .b(fc150), .c_in(fs166), .s(fs169), .c_out(fc169));

	logic fs170, fc170;
	FA fa170 (.a(fs167), .b(fc151), .c_in(fs168), .s(fs170), .c_out(fc170));

	logic fs171, fc171;
	FA fa171 (.a(fc152), .b(fs169), .c_in(fs170), .s(fs171), .c_out(fc171));

	logic hs21, hc21;
	HA ha21 (.a(in_0_21), .b(in_1_20), .s(hs21), .c_out(hc21));

	logic fs172, fc172;
	FA fa172 (.a(in_2_19), .b(in_3_18), .c_in(in_4_17), .s(fs172), .c_out(fc172));

	logic fs173, fc173;
	FA fa173 (.a(in_5_16), .b(in_6_15), .c_in(in_7_14), .s(fs173), .c_out(fc173));

	logic fs174, fc174;
	FA fa174 (.a(in_8_13), .b(in_9_12), .c_in(in_10_11), .s(fs174), .c_out(fc174));

	logic fs175, fc175;
	FA fa175 (.a(in_11_10), .b(in_12_9), .c_in(in_13_8), .s(fs175), .c_out(fc175));

	logic fs176, fc176;
	FA fa176 (.a(in_14_7), .b(in_15_6), .c_in(in_16_5), .s(fs176), .c_out(fc176));

	logic fs177, fc177;
	FA fa177 (.a(in_17_4), .b(in_18_3), .c_in(in_19_2), .s(fs177), .c_out(fc177));

	logic fs178, fc178;
	FA fa178 (.a(in_20_1), .b(in_21_0), .c_in(hc20), .s(fs178), .c_out(fc178));

	logic fs179, fc179;
	FA fa179 (.a(hs21), .b(fc154), .c_in(fc155), .s(fs179), .c_out(fc179));

	logic fs180, fc180;
	FA fa180 (.a(fc156), .b(fc157), .c_in(fc158), .s(fs180), .c_out(fc180));

	logic fs181, fc181;
	FA fa181 (.a(fc159), .b(fc160), .c_in(fs172), .s(fs181), .c_out(fc181));

	logic fs182, fc182;
	FA fa182 (.a(fs173), .b(fs174), .c_in(fs175), .s(fs182), .c_out(fc182));

	logic fs183, fc183;
	FA fa183 (.a(fs176), .b(fs177), .c_in(fs178), .s(fs183), .c_out(fc183));

	logic fs184, fc184;
	FA fa184 (.a(fc161), .b(fc162), .c_in(fc163), .s(fs184), .c_out(fc184));

	logic fs185, fc185;
	FA fa185 (.a(fc164), .b(fs179), .c_in(fs180), .s(fs185), .c_out(fc185));

	logic fs186, fc186;
	FA fa186 (.a(fc165), .b(fs181), .c_in(fs182), .s(fs186), .c_out(fc186));

	logic fs187, fc187;
	FA fa187 (.a(fs183), .b(fc166), .c_in(fc167), .s(fs187), .c_out(fc187));

	logic fs188, fc188;
	FA fa188 (.a(fs184), .b(fc168), .c_in(fs185), .s(fs188), .c_out(fc188));

	logic fs189, fc189;
	FA fa189 (.a(fs186), .b(fc169), .c_in(fs187), .s(fs189), .c_out(fc189));

	logic fs190, fc190;
	FA fa190 (.a(fc170), .b(fs188), .c_in(fs189), .s(fs190), .c_out(fc190));

	logic hs22, hc22;
	HA ha22 (.a(in_0_22), .b(in_1_21), .s(hs22), .c_out(hc22));

	logic fs191, fc191;
	FA fa191 (.a(in_2_20), .b(in_3_19), .c_in(in_4_18), .s(fs191), .c_out(fc191));

	logic fs192, fc192;
	FA fa192 (.a(in_5_17), .b(in_6_16), .c_in(in_7_15), .s(fs192), .c_out(fc192));

	logic fs193, fc193;
	FA fa193 (.a(in_8_14), .b(in_9_13), .c_in(in_10_12), .s(fs193), .c_out(fc193));

	logic fs194, fc194;
	FA fa194 (.a(in_11_11), .b(in_12_10), .c_in(in_13_9), .s(fs194), .c_out(fc194));

	logic fs195, fc195;
	FA fa195 (.a(in_14_8), .b(in_15_7), .c_in(in_16_6), .s(fs195), .c_out(fc195));

	logic fs196, fc196;
	FA fa196 (.a(in_17_5), .b(in_18_4), .c_in(in_19_3), .s(fs196), .c_out(fc196));

	logic fs197, fc197;
	FA fa197 (.a(in_20_2), .b(in_21_1), .c_in(in_22_0), .s(fs197), .c_out(fc197));

	logic fs198, fc198;
	FA fa198 (.a(hc21), .b(hs22), .c_in(fc172), .s(fs198), .c_out(fc198));

	logic fs199, fc199;
	FA fa199 (.a(fc173), .b(fc174), .c_in(fc175), .s(fs199), .c_out(fc199));

	logic fs200, fc200;
	FA fa200 (.a(fc176), .b(fc177), .c_in(fc178), .s(fs200), .c_out(fc200));

	logic fs201, fc201;
	FA fa201 (.a(fs191), .b(fs192), .c_in(fs193), .s(fs201), .c_out(fc201));

	logic fs202, fc202;
	FA fa202 (.a(fs194), .b(fs195), .c_in(fs196), .s(fs202), .c_out(fc202));

	logic fs203, fc203;
	FA fa203 (.a(fs197), .b(fc179), .c_in(fc180), .s(fs203), .c_out(fc203));

	logic fs204, fc204;
	FA fa204 (.a(fs198), .b(fc181), .c_in(fc182), .s(fs204), .c_out(fc204));

	logic fs205, fc205;
	FA fa205 (.a(fc183), .b(fs199), .c_in(fs200), .s(fs205), .c_out(fc205));

	logic fs206, fc206;
	FA fa206 (.a(fc184), .b(fs201), .c_in(fs202), .s(fs206), .c_out(fc206));

	logic fs207, fc207;
	FA fa207 (.a(fc185), .b(fs203), .c_in(fc186), .s(fs207), .c_out(fc207));

	logic fs208, fc208;
	FA fa208 (.a(fs204), .b(fs205), .c_in(fc187), .s(fs208), .c_out(fc208));

	logic fs209, fc209;
	FA fa209 (.a(fs206), .b(fc188), .c_in(fs207), .s(fs209), .c_out(fc209));

	logic fs210, fc210;
	FA fa210 (.a(fs208), .b(fc189), .c_in(fs209), .s(fs210), .c_out(fc210));

	logic hs23, hc23;
	HA ha23 (.a(in_0_23), .b(in_1_22), .s(hs23), .c_out(hc23));

	logic fs211, fc211;
	FA fa211 (.a(in_2_21), .b(in_3_20), .c_in(in_4_19), .s(fs211), .c_out(fc211));

	logic fs212, fc212;
	FA fa212 (.a(in_5_18), .b(in_6_17), .c_in(in_7_16), .s(fs212), .c_out(fc212));

	logic fs213, fc213;
	FA fa213 (.a(in_8_15), .b(in_9_14), .c_in(in_10_13), .s(fs213), .c_out(fc213));

	logic fs214, fc214;
	FA fa214 (.a(in_11_12), .b(in_12_11), .c_in(in_13_10), .s(fs214), .c_out(fc214));

	logic fs215, fc215;
	FA fa215 (.a(in_14_9), .b(in_15_8), .c_in(in_16_7), .s(fs215), .c_out(fc215));

	logic fs216, fc216;
	FA fa216 (.a(in_17_6), .b(in_18_5), .c_in(in_19_4), .s(fs216), .c_out(fc216));

	logic fs217, fc217;
	FA fa217 (.a(in_20_3), .b(in_21_2), .c_in(in_22_1), .s(fs217), .c_out(fc217));

	logic fs218, fc218;
	FA fa218 (.a(in_23_0), .b(hc22), .c_in(hs23), .s(fs218), .c_out(fc218));

	logic fs219, fc219;
	FA fa219 (.a(fc191), .b(fc192), .c_in(fc193), .s(fs219), .c_out(fc219));

	logic fs220, fc220;
	FA fa220 (.a(fc194), .b(fc195), .c_in(fc196), .s(fs220), .c_out(fc220));

	logic fs221, fc221;
	FA fa221 (.a(fc197), .b(fc198), .c_in(fs211), .s(fs221), .c_out(fc221));

	logic fs222, fc222;
	FA fa222 (.a(fs212), .b(fs213), .c_in(fs214), .s(fs222), .c_out(fc222));

	logic fs223, fc223;
	FA fa223 (.a(fs215), .b(fs216), .c_in(fs217), .s(fs223), .c_out(fc223));

	logic fs224, fc224;
	FA fa224 (.a(fs218), .b(fc199), .c_in(fc200), .s(fs224), .c_out(fc224));

	logic fs225, fc225;
	FA fa225 (.a(fc201), .b(fc202), .c_in(fs219), .s(fs225), .c_out(fc225));

	logic fs226, fc226;
	FA fa226 (.a(fs220), .b(fc203), .c_in(fs221), .s(fs226), .c_out(fc226));

	logic fs227, fc227;
	FA fa227 (.a(fs222), .b(fs223), .c_in(fc204), .s(fs227), .c_out(fc227));

	logic fs228, fc228;
	FA fa228 (.a(fc205), .b(fs224), .c_in(fc206), .s(fs228), .c_out(fc228));

	logic fs229, fc229;
	FA fa229 (.a(fs225), .b(fc207), .c_in(fs226), .s(fs229), .c_out(fc229));

	logic fs230, fc230;
	FA fa230 (.a(fs227), .b(fc208), .c_in(fs228), .s(fs230), .c_out(fc230));

	logic fs231, fc231;
	FA fa231 (.a(fc209), .b(fs229), .c_in(fs230), .s(fs231), .c_out(fc231));

	logic hs24, hc24;
	HA ha24 (.a(in_0_24), .b(in_1_23), .s(hs24), .c_out(hc24));

	logic fs232, fc232;
	FA fa232 (.a(in_2_22), .b(in_3_21), .c_in(in_4_20), .s(fs232), .c_out(fc232));

	logic fs233, fc233;
	FA fa233 (.a(in_5_19), .b(in_6_18), .c_in(in_7_17), .s(fs233), .c_out(fc233));

	logic fs234, fc234;
	FA fa234 (.a(in_8_16), .b(in_9_15), .c_in(in_10_14), .s(fs234), .c_out(fc234));

	logic fs235, fc235;
	FA fa235 (.a(in_11_13), .b(in_12_12), .c_in(in_13_11), .s(fs235), .c_out(fc235));

	logic fs236, fc236;
	FA fa236 (.a(in_14_10), .b(in_15_9), .c_in(in_16_8), .s(fs236), .c_out(fc236));

	logic fs237, fc237;
	FA fa237 (.a(in_17_7), .b(in_18_6), .c_in(in_19_5), .s(fs237), .c_out(fc237));

	logic fs238, fc238;
	FA fa238 (.a(in_20_4), .b(in_21_3), .c_in(in_22_2), .s(fs238), .c_out(fc238));

	logic fs239, fc239;
	FA fa239 (.a(in_23_1), .b(in_24_0), .c_in(hc23), .s(fs239), .c_out(fc239));

	logic fs240, fc240;
	FA fa240 (.a(hs24), .b(fc211), .c_in(fc212), .s(fs240), .c_out(fc240));

	logic fs241, fc241;
	FA fa241 (.a(fc213), .b(fc214), .c_in(fc215), .s(fs241), .c_out(fc241));

	logic fs242, fc242;
	FA fa242 (.a(fc216), .b(fc217), .c_in(fc218), .s(fs242), .c_out(fc242));

	logic fs243, fc243;
	FA fa243 (.a(fs232), .b(fs233), .c_in(fs234), .s(fs243), .c_out(fc243));

	logic fs244, fc244;
	FA fa244 (.a(fs235), .b(fs236), .c_in(fs237), .s(fs244), .c_out(fc244));

	logic fs245, fc245;
	FA fa245 (.a(fs238), .b(fs239), .c_in(fc219), .s(fs245), .c_out(fc245));

	logic fs246, fc246;
	FA fa246 (.a(fc220), .b(fc221), .c_in(fc222), .s(fs246), .c_out(fc246));

	logic fs247, fc247;
	FA fa247 (.a(fc223), .b(fs240), .c_in(fs241), .s(fs247), .c_out(fc247));

	logic fs248, fc248;
	FA fa248 (.a(fs242), .b(fc224), .c_in(fs243), .s(fs248), .c_out(fc248));

	logic fs249, fc249;
	FA fa249 (.a(fs244), .b(fs245), .c_in(fc225), .s(fs249), .c_out(fc249));

	logic fs250, fc250;
	FA fa250 (.a(fc226), .b(fc227), .c_in(fs246), .s(fs250), .c_out(fc250));

	logic fs251, fc251;
	FA fa251 (.a(fs247), .b(fc228), .c_in(fs248), .s(fs251), .c_out(fc251));

	logic fs252, fc252;
	FA fa252 (.a(fs249), .b(fc229), .c_in(fs250), .s(fs252), .c_out(fc252));

	logic fs253, fc253;
	FA fa253 (.a(fc230), .b(fs251), .c_in(fs252), .s(fs253), .c_out(fc253));

	logic hs25, hc25;
	HA ha25 (.a(in_0_25), .b(in_1_24), .s(hs25), .c_out(hc25));

	logic fs254, fc254;
	FA fa254 (.a(in_2_23), .b(in_3_22), .c_in(in_4_21), .s(fs254), .c_out(fc254));

	logic fs255, fc255;
	FA fa255 (.a(in_5_20), .b(in_6_19), .c_in(in_7_18), .s(fs255), .c_out(fc255));

	logic fs256, fc256;
	FA fa256 (.a(in_8_17), .b(in_9_16), .c_in(in_10_15), .s(fs256), .c_out(fc256));

	logic fs257, fc257;
	FA fa257 (.a(in_11_14), .b(in_12_13), .c_in(in_13_12), .s(fs257), .c_out(fc257));

	logic fs258, fc258;
	FA fa258 (.a(in_14_11), .b(in_15_10), .c_in(in_16_9), .s(fs258), .c_out(fc258));

	logic fs259, fc259;
	FA fa259 (.a(in_17_8), .b(in_18_7), .c_in(in_19_6), .s(fs259), .c_out(fc259));

	logic fs260, fc260;
	FA fa260 (.a(in_20_5), .b(in_21_4), .c_in(in_22_3), .s(fs260), .c_out(fc260));

	logic fs261, fc261;
	FA fa261 (.a(in_23_2), .b(in_24_1), .c_in(in_25_0), .s(fs261), .c_out(fc261));

	logic fs262, fc262;
	FA fa262 (.a(hc24), .b(hs25), .c_in(fc232), .s(fs262), .c_out(fc262));

	logic fs263, fc263;
	FA fa263 (.a(fc233), .b(fc234), .c_in(fc235), .s(fs263), .c_out(fc263));

	logic fs264, fc264;
	FA fa264 (.a(fc236), .b(fc237), .c_in(fc238), .s(fs264), .c_out(fc264));

	logic fs265, fc265;
	FA fa265 (.a(fc239), .b(fs254), .c_in(fs255), .s(fs265), .c_out(fc265));

	logic fs266, fc266;
	FA fa266 (.a(fs256), .b(fs257), .c_in(fs258), .s(fs266), .c_out(fc266));

	logic fs267, fc267;
	FA fa267 (.a(fs259), .b(fs260), .c_in(fs261), .s(fs267), .c_out(fc267));

	logic fs268, fc268;
	FA fa268 (.a(fc240), .b(fc241), .c_in(fc242), .s(fs268), .c_out(fc268));

	logic fs269, fc269;
	FA fa269 (.a(fs262), .b(fc243), .c_in(fc244), .s(fs269), .c_out(fc269));

	logic fs270, fc270;
	FA fa270 (.a(fc245), .b(fs263), .c_in(fs264), .s(fs270), .c_out(fc270));

	logic fs271, fc271;
	FA fa271 (.a(fs265), .b(fs266), .c_in(fs267), .s(fs271), .c_out(fc271));

	logic fs272, fc272;
	FA fa272 (.a(fc246), .b(fc247), .c_in(fs268), .s(fs272), .c_out(fc272));

	logic fs273, fc273;
	FA fa273 (.a(fc248), .b(fc249), .c_in(fs269), .s(fs273), .c_out(fc273));

	logic fs274, fc274;
	FA fa274 (.a(fs270), .b(fs271), .c_in(fc250), .s(fs274), .c_out(fc274));

	logic fs275, fc275;
	FA fa275 (.a(fs272), .b(fc251), .c_in(fs273), .s(fs275), .c_out(fc275));

	logic fs276, fc276;
	FA fa276 (.a(fs274), .b(fc252), .c_in(fs275), .s(fs276), .c_out(fc276));

	logic hs26, hc26;
	HA ha26 (.a(in_0_26), .b(in_1_25), .s(hs26), .c_out(hc26));

	logic fs277, fc277;
	FA fa277 (.a(in_2_24), .b(in_3_23), .c_in(in_4_22), .s(fs277), .c_out(fc277));

	logic fs278, fc278;
	FA fa278 (.a(in_5_21), .b(in_6_20), .c_in(in_7_19), .s(fs278), .c_out(fc278));

	logic fs279, fc279;
	FA fa279 (.a(in_8_18), .b(in_9_17), .c_in(in_10_16), .s(fs279), .c_out(fc279));

	logic fs280, fc280;
	FA fa280 (.a(in_11_15), .b(in_12_14), .c_in(in_13_13), .s(fs280), .c_out(fc280));

	logic fs281, fc281;
	FA fa281 (.a(in_14_12), .b(in_15_11), .c_in(in_16_10), .s(fs281), .c_out(fc281));

	logic fs282, fc282;
	FA fa282 (.a(in_17_9), .b(in_18_8), .c_in(in_19_7), .s(fs282), .c_out(fc282));

	logic fs283, fc283;
	FA fa283 (.a(in_20_6), .b(in_21_5), .c_in(in_22_4), .s(fs283), .c_out(fc283));

	logic fs284, fc284;
	FA fa284 (.a(in_23_3), .b(in_24_2), .c_in(in_25_1), .s(fs284), .c_out(fc284));

	logic fs285, fc285;
	FA fa285 (.a(in_26_0), .b(hc25), .c_in(hs26), .s(fs285), .c_out(fc285));

	logic fs286, fc286;
	FA fa286 (.a(fc254), .b(fc255), .c_in(fc256), .s(fs286), .c_out(fc286));

	logic fs287, fc287;
	FA fa287 (.a(fc257), .b(fc258), .c_in(fc259), .s(fs287), .c_out(fc287));

	logic fs288, fc288;
	FA fa288 (.a(fc260), .b(fc261), .c_in(fc262), .s(fs288), .c_out(fc288));

	logic fs289, fc289;
	FA fa289 (.a(fs277), .b(fs278), .c_in(fs279), .s(fs289), .c_out(fc289));

	logic fs290, fc290;
	FA fa290 (.a(fs280), .b(fs281), .c_in(fs282), .s(fs290), .c_out(fc290));

	logic fs291, fc291;
	FA fa291 (.a(fs283), .b(fs284), .c_in(fs285), .s(fs291), .c_out(fc291));

	logic fs292, fc292;
	FA fa292 (.a(fc263), .b(fc264), .c_in(fc265), .s(fs292), .c_out(fc292));

	logic fs293, fc293;
	FA fa293 (.a(fc266), .b(fc267), .c_in(fs286), .s(fs293), .c_out(fc293));

	logic fs294, fc294;
	FA fa294 (.a(fs287), .b(fs288), .c_in(fc268), .s(fs294), .c_out(fc294));

	logic fs295, fc295;
	FA fa295 (.a(fs289), .b(fs290), .c_in(fs291), .s(fs295), .c_out(fc295));

	logic fs296, fc296;
	FA fa296 (.a(fc269), .b(fc270), .c_in(fs292), .s(fs296), .c_out(fc296));

	logic fs297, fc297;
	FA fa297 (.a(fc271), .b(fs293), .c_in(fs294), .s(fs297), .c_out(fc297));

	logic fs298, fc298;
	FA fa298 (.a(fc272), .b(fs295), .c_in(fc273), .s(fs298), .c_out(fc298));

	logic fs299, fc299;
	FA fa299 (.a(fs296), .b(fc274), .c_in(fs297), .s(fs299), .c_out(fc299));

	logic fs300, fc300;
	FA fa300 (.a(fs298), .b(fc275), .c_in(fs299), .s(fs300), .c_out(fc300));

	logic hs27, hc27;
	HA ha27 (.a(in_0_27), .b(in_1_26), .s(hs27), .c_out(hc27));

	logic fs301, fc301;
	FA fa301 (.a(in_2_25), .b(in_3_24), .c_in(in_4_23), .s(fs301), .c_out(fc301));

	logic fs302, fc302;
	FA fa302 (.a(in_5_22), .b(in_6_21), .c_in(in_7_20), .s(fs302), .c_out(fc302));

	logic fs303, fc303;
	FA fa303 (.a(in_8_19), .b(in_9_18), .c_in(in_10_17), .s(fs303), .c_out(fc303));

	logic fs304, fc304;
	FA fa304 (.a(in_11_16), .b(in_12_15), .c_in(in_13_14), .s(fs304), .c_out(fc304));

	logic fs305, fc305;
	FA fa305 (.a(in_14_13), .b(in_15_12), .c_in(in_16_11), .s(fs305), .c_out(fc305));

	logic fs306, fc306;
	FA fa306 (.a(in_17_10), .b(in_18_9), .c_in(in_19_8), .s(fs306), .c_out(fc306));

	logic fs307, fc307;
	FA fa307 (.a(in_20_7), .b(in_21_6), .c_in(in_22_5), .s(fs307), .c_out(fc307));

	logic fs308, fc308;
	FA fa308 (.a(in_23_4), .b(in_24_3), .c_in(in_25_2), .s(fs308), .c_out(fc308));

	logic fs309, fc309;
	FA fa309 (.a(in_26_1), .b(in_27_0), .c_in(hc26), .s(fs309), .c_out(fc309));

	logic fs310, fc310;
	FA fa310 (.a(hs27), .b(fc277), .c_in(fc278), .s(fs310), .c_out(fc310));

	logic fs311, fc311;
	FA fa311 (.a(fc279), .b(fc280), .c_in(fc281), .s(fs311), .c_out(fc311));

	logic fs312, fc312;
	FA fa312 (.a(fc282), .b(fc283), .c_in(fc284), .s(fs312), .c_out(fc312));

	logic fs313, fc313;
	FA fa313 (.a(fc285), .b(fs301), .c_in(fs302), .s(fs313), .c_out(fc313));

	logic fs314, fc314;
	FA fa314 (.a(fs303), .b(fs304), .c_in(fs305), .s(fs314), .c_out(fc314));

	logic fs315, fc315;
	FA fa315 (.a(fs306), .b(fs307), .c_in(fs308), .s(fs315), .c_out(fc315));

	logic fs316, fc316;
	FA fa316 (.a(fs309), .b(fc286), .c_in(fc287), .s(fs316), .c_out(fc316));

	logic fs317, fc317;
	FA fa317 (.a(fc288), .b(fc289), .c_in(fc290), .s(fs317), .c_out(fc317));

	logic fs318, fc318;
	FA fa318 (.a(fc291), .b(fs310), .c_in(fs311), .s(fs318), .c_out(fc318));

	logic fs319, fc319;
	FA fa319 (.a(fs312), .b(fc292), .c_in(fs313), .s(fs319), .c_out(fc319));

	logic fs320, fc320;
	FA fa320 (.a(fs314), .b(fs315), .c_in(fc293), .s(fs320), .c_out(fc320));

	logic fs321, fc321;
	FA fa321 (.a(fc294), .b(fs316), .c_in(fc295), .s(fs321), .c_out(fc321));

	logic fs322, fc322;
	FA fa322 (.a(fs317), .b(fs318), .c_in(fc296), .s(fs322), .c_out(fc322));

	logic fs323, fc323;
	FA fa323 (.a(fs319), .b(fs320), .c_in(fc297), .s(fs323), .c_out(fc323));

	logic fs324, fc324;
	FA fa324 (.a(fs321), .b(fc298), .c_in(fs322), .s(fs324), .c_out(fc324));

	logic fs325, fc325;
	FA fa325 (.a(fs323), .b(fc299), .c_in(fs324), .s(fs325), .c_out(fc325));

	logic hs28, hc28;
	HA ha28 (.a(in_0_28), .b(in_1_27), .s(hs28), .c_out(hc28));

	logic fs326, fc326;
	FA fa326 (.a(in_2_26), .b(in_3_25), .c_in(in_4_24), .s(fs326), .c_out(fc326));

	logic fs327, fc327;
	FA fa327 (.a(in_5_23), .b(in_6_22), .c_in(in_7_21), .s(fs327), .c_out(fc327));

	logic fs328, fc328;
	FA fa328 (.a(in_8_20), .b(in_9_19), .c_in(in_10_18), .s(fs328), .c_out(fc328));

	logic fs329, fc329;
	FA fa329 (.a(in_11_17), .b(in_12_16), .c_in(in_13_15), .s(fs329), .c_out(fc329));

	logic fs330, fc330;
	FA fa330 (.a(in_14_14), .b(in_15_13), .c_in(in_16_12), .s(fs330), .c_out(fc330));

	logic fs331, fc331;
	FA fa331 (.a(in_17_11), .b(in_18_10), .c_in(in_19_9), .s(fs331), .c_out(fc331));

	logic fs332, fc332;
	FA fa332 (.a(in_20_8), .b(in_21_7), .c_in(in_22_6), .s(fs332), .c_out(fc332));

	logic fs333, fc333;
	FA fa333 (.a(in_23_5), .b(in_24_4), .c_in(in_25_3), .s(fs333), .c_out(fc333));

	logic fs334, fc334;
	FA fa334 (.a(in_26_2), .b(in_27_1), .c_in(in_28_0), .s(fs334), .c_out(fc334));

	logic fs335, fc335;
	FA fa335 (.a(hc27), .b(hs28), .c_in(fc301), .s(fs335), .c_out(fc335));

	logic fs336, fc336;
	FA fa336 (.a(fc302), .b(fc303), .c_in(fc304), .s(fs336), .c_out(fc336));

	logic fs337, fc337;
	FA fa337 (.a(fc305), .b(fc306), .c_in(fc307), .s(fs337), .c_out(fc337));

	logic fs338, fc338;
	FA fa338 (.a(fc308), .b(fc309), .c_in(fs326), .s(fs338), .c_out(fc338));

	logic fs339, fc339;
	FA fa339 (.a(fs327), .b(fs328), .c_in(fs329), .s(fs339), .c_out(fc339));

	logic fs340, fc340;
	FA fa340 (.a(fs330), .b(fs331), .c_in(fs332), .s(fs340), .c_out(fc340));

	logic fs341, fc341;
	FA fa341 (.a(fs333), .b(fs334), .c_in(fc310), .s(fs341), .c_out(fc341));

	logic fs342, fc342;
	FA fa342 (.a(fc311), .b(fc312), .c_in(fs335), .s(fs342), .c_out(fc342));

	logic fs343, fc343;
	FA fa343 (.a(fc313), .b(fc314), .c_in(fc315), .s(fs343), .c_out(fc343));

	logic fs344, fc344;
	FA fa344 (.a(fs336), .b(fs337), .c_in(fs338), .s(fs344), .c_out(fc344));

	logic fs345, fc345;
	FA fa345 (.a(fc316), .b(fs339), .c_in(fs340), .s(fs345), .c_out(fc345));

	logic fs346, fc346;
	FA fa346 (.a(fs341), .b(fc317), .c_in(fc318), .s(fs346), .c_out(fc346));

	logic fs347, fc347;
	FA fa347 (.a(fs342), .b(fc319), .c_in(fc320), .s(fs347), .c_out(fc347));

	logic fs348, fc348;
	FA fa348 (.a(fs343), .b(fs344), .c_in(fc321), .s(fs348), .c_out(fc348));

	logic fs349, fc349;
	FA fa349 (.a(fs345), .b(fc322), .c_in(fs346), .s(fs349), .c_out(fc349));

	logic fs350, fc350;
	FA fa350 (.a(fc323), .b(fs347), .c_in(fs348), .s(fs350), .c_out(fc350));

	logic fs351, fc351;
	FA fa351 (.a(fc324), .b(fs349), .c_in(fs350), .s(fs351), .c_out(fc351));

	logic hs29, hc29;
	HA ha29 (.a(in_0_29), .b(in_1_28), .s(hs29), .c_out(hc29));

	logic fs352, fc352;
	FA fa352 (.a(in_2_27), .b(in_3_26), .c_in(in_4_25), .s(fs352), .c_out(fc352));

	logic fs353, fc353;
	FA fa353 (.a(in_5_24), .b(in_6_23), .c_in(in_7_22), .s(fs353), .c_out(fc353));

	logic fs354, fc354;
	FA fa354 (.a(in_8_21), .b(in_9_20), .c_in(in_10_19), .s(fs354), .c_out(fc354));

	logic fs355, fc355;
	FA fa355 (.a(in_11_18), .b(in_12_17), .c_in(in_13_16), .s(fs355), .c_out(fc355));

	logic fs356, fc356;
	FA fa356 (.a(in_14_15), .b(in_15_14), .c_in(in_16_13), .s(fs356), .c_out(fc356));

	logic fs357, fc357;
	FA fa357 (.a(in_17_12), .b(in_18_11), .c_in(in_19_10), .s(fs357), .c_out(fc357));

	logic fs358, fc358;
	FA fa358 (.a(in_20_9), .b(in_21_8), .c_in(in_22_7), .s(fs358), .c_out(fc358));

	logic fs359, fc359;
	FA fa359 (.a(in_23_6), .b(in_24_5), .c_in(in_25_4), .s(fs359), .c_out(fc359));

	logic fs360, fc360;
	FA fa360 (.a(in_26_3), .b(in_27_2), .c_in(in_28_1), .s(fs360), .c_out(fc360));

	logic fs361, fc361;
	FA fa361 (.a(in_29_0), .b(hc28), .c_in(hs29), .s(fs361), .c_out(fc361));

	logic fs362, fc362;
	FA fa362 (.a(fc326), .b(fc327), .c_in(fc328), .s(fs362), .c_out(fc362));

	logic fs363, fc363;
	FA fa363 (.a(fc329), .b(fc330), .c_in(fc331), .s(fs363), .c_out(fc363));

	logic fs364, fc364;
	FA fa364 (.a(fc332), .b(fc333), .c_in(fc334), .s(fs364), .c_out(fc364));

	logic fs365, fc365;
	FA fa365 (.a(fc335), .b(fs352), .c_in(fs353), .s(fs365), .c_out(fc365));

	logic fs366, fc366;
	FA fa366 (.a(fs354), .b(fs355), .c_in(fs356), .s(fs366), .c_out(fc366));

	logic fs367, fc367;
	FA fa367 (.a(fs357), .b(fs358), .c_in(fs359), .s(fs367), .c_out(fc367));

	logic fs368, fc368;
	FA fa368 (.a(fs360), .b(fs361), .c_in(fc336), .s(fs368), .c_out(fc368));

	logic fs369, fc369;
	FA fa369 (.a(fc337), .b(fc338), .c_in(fc339), .s(fs369), .c_out(fc369));

	logic fs370, fc370;
	FA fa370 (.a(fc340), .b(fc341), .c_in(fs362), .s(fs370), .c_out(fc370));

	logic fs371, fc371;
	FA fa371 (.a(fs363), .b(fs364), .c_in(fc342), .s(fs371), .c_out(fc371));

	logic fs372, fc372;
	FA fa372 (.a(fs365), .b(fs366), .c_in(fs367), .s(fs372), .c_out(fc372));

	logic fs373, fc373;
	FA fa373 (.a(fs368), .b(fc343), .c_in(fc344), .s(fs373), .c_out(fc373));

	logic fs374, fc374;
	FA fa374 (.a(fs369), .b(fc345), .c_in(fs370), .s(fs374), .c_out(fc374));

	logic fs375, fc375;
	FA fa375 (.a(fs371), .b(fc346), .c_in(fs372), .s(fs375), .c_out(fc375));

	logic fs376, fc376;
	FA fa376 (.a(fc347), .b(fc348), .c_in(fs373), .s(fs376), .c_out(fc376));

	logic fs377, fc377;
	FA fa377 (.a(fs374), .b(fc349), .c_in(fs375), .s(fs377), .c_out(fc377));

	logic fs378, fc378;
	FA fa378 (.a(fc350), .b(fs376), .c_in(fs377), .s(fs378), .c_out(fc378));

	logic hs30, hc30;
	HA ha30 (.a(in_0_30), .b(in_1_29), .s(hs30), .c_out(hc30));

	logic fs379, fc379;
	FA fa379 (.a(in_2_28), .b(in_3_27), .c_in(in_4_26), .s(fs379), .c_out(fc379));

	logic fs380, fc380;
	FA fa380 (.a(in_5_25), .b(in_6_24), .c_in(in_7_23), .s(fs380), .c_out(fc380));

	logic fs381, fc381;
	FA fa381 (.a(in_8_22), .b(in_9_21), .c_in(in_10_20), .s(fs381), .c_out(fc381));

	logic fs382, fc382;
	FA fa382 (.a(in_11_19), .b(in_12_18), .c_in(in_13_17), .s(fs382), .c_out(fc382));

	logic fs383, fc383;
	FA fa383 (.a(in_14_16), .b(in_15_15), .c_in(in_16_14), .s(fs383), .c_out(fc383));

	logic fs384, fc384;
	FA fa384 (.a(in_17_13), .b(in_18_12), .c_in(in_19_11), .s(fs384), .c_out(fc384));

	logic fs385, fc385;
	FA fa385 (.a(in_20_10), .b(in_21_9), .c_in(in_22_8), .s(fs385), .c_out(fc385));

	logic fs386, fc386;
	FA fa386 (.a(in_23_7), .b(in_24_6), .c_in(in_25_5), .s(fs386), .c_out(fc386));

	logic fs387, fc387;
	FA fa387 (.a(in_26_4), .b(in_27_3), .c_in(in_28_2), .s(fs387), .c_out(fc387));

	logic fs388, fc388;
	FA fa388 (.a(in_29_1), .b(in_30_0), .c_in(hc29), .s(fs388), .c_out(fc388));

	logic fs389, fc389;
	FA fa389 (.a(hs30), .b(fc352), .c_in(fc353), .s(fs389), .c_out(fc389));

	logic fs390, fc390;
	FA fa390 (.a(fc354), .b(fc355), .c_in(fc356), .s(fs390), .c_out(fc390));

	logic fs391, fc391;
	FA fa391 (.a(fc357), .b(fc358), .c_in(fc359), .s(fs391), .c_out(fc391));

	logic fs392, fc392;
	FA fa392 (.a(fc360), .b(fc361), .c_in(fs379), .s(fs392), .c_out(fc392));

	logic fs393, fc393;
	FA fa393 (.a(fs380), .b(fs381), .c_in(fs382), .s(fs393), .c_out(fc393));

	logic fs394, fc394;
	FA fa394 (.a(fs383), .b(fs384), .c_in(fs385), .s(fs394), .c_out(fc394));

	logic fs395, fc395;
	FA fa395 (.a(fs386), .b(fs387), .c_in(fs388), .s(fs395), .c_out(fc395));

	logic fs396, fc396;
	FA fa396 (.a(fc362), .b(fc363), .c_in(fc364), .s(fs396), .c_out(fc396));

	logic fs397, fc397;
	FA fa397 (.a(fc365), .b(fc366), .c_in(fc367), .s(fs397), .c_out(fc397));

	logic fs398, fc398;
	FA fa398 (.a(fs389), .b(fs390), .c_in(fs391), .s(fs398), .c_out(fc398));

	logic fs399, fc399;
	FA fa399 (.a(fc368), .b(fs392), .c_in(fc369), .s(fs399), .c_out(fc399));

	logic fs400, fc400;
	FA fa400 (.a(fs393), .b(fs394), .c_in(fs395), .s(fs400), .c_out(fc400));

	logic fs401, fc401;
	FA fa401 (.a(fc370), .b(fc371), .c_in(fs396), .s(fs401), .c_out(fc401));

	logic fs402, fc402;
	FA fa402 (.a(fc372), .b(fs397), .c_in(fs398), .s(fs402), .c_out(fc402));

	logic fs403, fc403;
	FA fa403 (.a(fs399), .b(fc373), .c_in(fs400), .s(fs403), .c_out(fc403));

	logic fs404, fc404;
	FA fa404 (.a(fc374), .b(fs401), .c_in(fc375), .s(fs404), .c_out(fc404));

	logic fs405, fc405;
	FA fa405 (.a(fs402), .b(fc376), .c_in(fs403), .s(fs405), .c_out(fc405));

	logic fs406, fc406;
	FA fa406 (.a(fs404), .b(fc377), .c_in(fs405), .s(fs406), .c_out(fc406));

	logic hs31, hc31;
	HA ha31 (.a(in_0_31), .b(in_1_30), .s(hs31), .c_out(hc31));

	logic fs407, fc407;
	FA fa407 (.a(in_2_29), .b(in_3_28), .c_in(in_4_27), .s(fs407), .c_out(fc407));

	logic fs408, fc408;
	FA fa408 (.a(in_5_26), .b(in_6_25), .c_in(in_7_24), .s(fs408), .c_out(fc408));

	logic fs409, fc409;
	FA fa409 (.a(in_8_23), .b(in_9_22), .c_in(in_10_21), .s(fs409), .c_out(fc409));

	logic fs410, fc410;
	FA fa410 (.a(in_11_20), .b(in_12_19), .c_in(in_13_18), .s(fs410), .c_out(fc410));

	logic fs411, fc411;
	FA fa411 (.a(in_14_17), .b(in_15_16), .c_in(in_16_15), .s(fs411), .c_out(fc411));

	logic fs412, fc412;
	FA fa412 (.a(in_17_14), .b(in_18_13), .c_in(in_19_12), .s(fs412), .c_out(fc412));

	logic fs413, fc413;
	FA fa413 (.a(in_20_11), .b(in_21_10), .c_in(in_22_9), .s(fs413), .c_out(fc413));

	logic fs414, fc414;
	FA fa414 (.a(in_23_8), .b(in_24_7), .c_in(in_25_6), .s(fs414), .c_out(fc414));

	logic fs415, fc415;
	FA fa415 (.a(in_26_5), .b(in_27_4), .c_in(in_28_3), .s(fs415), .c_out(fc415));

	logic fs416, fc416;
	FA fa416 (.a(in_29_2), .b(in_30_1), .c_in(in_31_0), .s(fs416), .c_out(fc416));

	logic fs417, fc417;
	FA fa417 (.a(hc30), .b(hs31), .c_in(fc379), .s(fs417), .c_out(fc417));

	logic fs418, fc418;
	FA fa418 (.a(fc380), .b(fc381), .c_in(fc382), .s(fs418), .c_out(fc418));

	logic fs419, fc419;
	FA fa419 (.a(fc383), .b(fc384), .c_in(fc385), .s(fs419), .c_out(fc419));

	logic fs420, fc420;
	FA fa420 (.a(fc386), .b(fc387), .c_in(fc388), .s(fs420), .c_out(fc420));

	logic fs421, fc421;
	FA fa421 (.a(fs407), .b(fs408), .c_in(fs409), .s(fs421), .c_out(fc421));

	logic fs422, fc422;
	FA fa422 (.a(fs410), .b(fs411), .c_in(fs412), .s(fs422), .c_out(fc422));

	logic fs423, fc423;
	FA fa423 (.a(fs413), .b(fs414), .c_in(fs415), .s(fs423), .c_out(fc423));

	logic fs424, fc424;
	FA fa424 (.a(fs416), .b(fc389), .c_in(fc390), .s(fs424), .c_out(fc424));

	logic fs425, fc425;
	FA fa425 (.a(fc391), .b(fs417), .c_in(fc392), .s(fs425), .c_out(fc425));

	logic fs426, fc426;
	FA fa426 (.a(fc393), .b(fc394), .c_in(fc395), .s(fs426), .c_out(fc426));

	logic fs427, fc427;
	FA fa427 (.a(fs418), .b(fs419), .c_in(fs420), .s(fs427), .c_out(fc427));

	logic fs428, fc428;
	FA fa428 (.a(fc396), .b(fs421), .c_in(fs422), .s(fs428), .c_out(fc428));

	logic fs429, fc429;
	FA fa429 (.a(fs423), .b(fc397), .c_in(fc398), .s(fs429), .c_out(fc429));

	logic fs430, fc430;
	FA fa430 (.a(fs424), .b(fs425), .c_in(fc399), .s(fs430), .c_out(fc430));

	logic fs431, fc431;
	FA fa431 (.a(fc400), .b(fs426), .c_in(fs427), .s(fs431), .c_out(fc431));

	logic fs432, fc432;
	FA fa432 (.a(fc401), .b(fs428), .c_in(fc402), .s(fs432), .c_out(fc432));

	logic fs433, fc433;
	FA fa433 (.a(fs429), .b(fs430), .c_in(fc403), .s(fs433), .c_out(fc433));

	logic fs434, fc434;
	FA fa434 (.a(fs431), .b(fc404), .c_in(fs432), .s(fs434), .c_out(fc434));

	logic fs435, fc435;
	FA fa435 (.a(fs433), .b(fc405), .c_in(fs434), .s(fs435), .c_out(fc435));

	logic hs32, hc32;
	HA ha32 (.a(in_1_31), .b(in_2_30), .s(hs32), .c_out(hc32));

	logic fs436, fc436;
	FA fa436 (.a(in_3_29), .b(in_4_28), .c_in(in_5_27), .s(fs436), .c_out(fc436));

	logic fs437, fc437;
	FA fa437 (.a(in_6_26), .b(in_7_25), .c_in(in_8_24), .s(fs437), .c_out(fc437));

	logic fs438, fc438;
	FA fa438 (.a(in_9_23), .b(in_10_22), .c_in(in_11_21), .s(fs438), .c_out(fc438));

	logic fs439, fc439;
	FA fa439 (.a(in_12_20), .b(in_13_19), .c_in(in_14_18), .s(fs439), .c_out(fc439));

	logic fs440, fc440;
	FA fa440 (.a(in_15_17), .b(in_16_16), .c_in(in_17_15), .s(fs440), .c_out(fc440));

	logic fs441, fc441;
	FA fa441 (.a(in_18_14), .b(in_19_13), .c_in(in_20_12), .s(fs441), .c_out(fc441));

	logic fs442, fc442;
	FA fa442 (.a(in_21_11), .b(in_22_10), .c_in(in_23_9), .s(fs442), .c_out(fc442));

	logic fs443, fc443;
	FA fa443 (.a(in_24_8), .b(in_25_7), .c_in(in_26_6), .s(fs443), .c_out(fc443));

	logic fs444, fc444;
	FA fa444 (.a(in_27_5), .b(in_28_4), .c_in(in_29_3), .s(fs444), .c_out(fc444));

	logic fs445, fc445;
	FA fa445 (.a(in_30_2), .b(in_31_1), .c_in(hc31), .s(fs445), .c_out(fc445));

	logic fs446, fc446;
	FA fa446 (.a(hs32), .b(fc407), .c_in(fc408), .s(fs446), .c_out(fc446));

	logic fs447, fc447;
	FA fa447 (.a(fc409), .b(fc410), .c_in(fc411), .s(fs447), .c_out(fc447));

	logic fs448, fc448;
	FA fa448 (.a(fc412), .b(fc413), .c_in(fc414), .s(fs448), .c_out(fc448));

	logic fs449, fc449;
	FA fa449 (.a(fc415), .b(fc416), .c_in(fc417), .s(fs449), .c_out(fc449));

	logic fs450, fc450;
	FA fa450 (.a(fs436), .b(fs437), .c_in(fs438), .s(fs450), .c_out(fc450));

	logic fs451, fc451;
	FA fa451 (.a(fs439), .b(fs440), .c_in(fs441), .s(fs451), .c_out(fc451));

	logic fs452, fc452;
	FA fa452 (.a(fs442), .b(fs443), .c_in(fs444), .s(fs452), .c_out(fc452));

	logic fs453, fc453;
	FA fa453 (.a(fs445), .b(fc418), .c_in(fc419), .s(fs453), .c_out(fc453));

	logic fs454, fc454;
	FA fa454 (.a(fc420), .b(fc421), .c_in(fc422), .s(fs454), .c_out(fc454));

	logic fs455, fc455;
	FA fa455 (.a(fc423), .b(fs446), .c_in(fs447), .s(fs455), .c_out(fc455));

	logic fs456, fc456;
	FA fa456 (.a(fs448), .b(fs449), .c_in(fc424), .s(fs456), .c_out(fc456));

	logic fs457, fc457;
	FA fa457 (.a(fc425), .b(fs450), .c_in(fs451), .s(fs457), .c_out(fc457));

	logic fs458, fc458;
	FA fa458 (.a(fs452), .b(fc426), .c_in(fc427), .s(fs458), .c_out(fc458));

	logic fs459, fc459;
	FA fa459 (.a(fs453), .b(fc428), .c_in(fs454), .s(fs459), .c_out(fc459));

	logic fs460, fc460;
	FA fa460 (.a(fs455), .b(fs456), .c_in(fc429), .s(fs460), .c_out(fc460));

	logic fs461, fc461;
	FA fa461 (.a(fc430), .b(fs457), .c_in(fc431), .s(fs461), .c_out(fc461));

	logic fs462, fc462;
	FA fa462 (.a(fs458), .b(fc432), .c_in(fs459), .s(fs462), .c_out(fc462));

	logic fs463, fc463;
	FA fa463 (.a(fs460), .b(fc433), .c_in(fs461), .s(fs463), .c_out(fc463));

	logic fs464, fc464;
	FA fa464 (.a(fc434), .b(fs462), .c_in(fs463), .s(fs464), .c_out(fc464));

	logic fs465, fc465;
	FA fa465 (.a(in_2_31), .b(in_3_30), .c_in(in_4_29), .s(fs465), .c_out(fc465));

	logic fs466, fc466;
	FA fa466 (.a(in_5_28), .b(in_6_27), .c_in(in_7_26), .s(fs466), .c_out(fc466));

	logic fs467, fc467;
	FA fa467 (.a(in_8_25), .b(in_9_24), .c_in(in_10_23), .s(fs467), .c_out(fc467));

	logic fs468, fc468;
	FA fa468 (.a(in_11_22), .b(in_12_21), .c_in(in_13_20), .s(fs468), .c_out(fc468));

	logic fs469, fc469;
	FA fa469 (.a(in_14_19), .b(in_15_18), .c_in(in_16_17), .s(fs469), .c_out(fc469));

	logic fs470, fc470;
	FA fa470 (.a(in_17_16), .b(in_18_15), .c_in(in_19_14), .s(fs470), .c_out(fc470));

	logic fs471, fc471;
	FA fa471 (.a(in_20_13), .b(in_21_12), .c_in(in_22_11), .s(fs471), .c_out(fc471));

	logic fs472, fc472;
	FA fa472 (.a(in_23_10), .b(in_24_9), .c_in(in_25_8), .s(fs472), .c_out(fc472));

	logic fs473, fc473;
	FA fa473 (.a(in_26_7), .b(in_27_6), .c_in(in_28_5), .s(fs473), .c_out(fc473));

	logic fs474, fc474;
	FA fa474 (.a(in_29_4), .b(in_30_3), .c_in(in_31_2), .s(fs474), .c_out(fc474));

	logic fs475, fc475;
	FA fa475 (.a(hc32), .b(fc436), .c_in(fc437), .s(fs475), .c_out(fc475));

	logic fs476, fc476;
	FA fa476 (.a(fc438), .b(fc439), .c_in(fc440), .s(fs476), .c_out(fc476));

	logic fs477, fc477;
	FA fa477 (.a(fc441), .b(fc442), .c_in(fc443), .s(fs477), .c_out(fc477));

	logic fs478, fc478;
	FA fa478 (.a(fc444), .b(fc445), .c_in(fs465), .s(fs478), .c_out(fc478));

	logic fs479, fc479;
	FA fa479 (.a(fs466), .b(fs467), .c_in(fs468), .s(fs479), .c_out(fc479));

	logic fs480, fc480;
	FA fa480 (.a(fs469), .b(fs470), .c_in(fs471), .s(fs480), .c_out(fc480));

	logic fs481, fc481;
	FA fa481 (.a(fs472), .b(fs473), .c_in(fs474), .s(fs481), .c_out(fc481));

	logic fs482, fc482;
	FA fa482 (.a(fc446), .b(fc447), .c_in(fc448), .s(fs482), .c_out(fc482));

	logic fs483, fc483;
	FA fa483 (.a(fc449), .b(fc450), .c_in(fc451), .s(fs483), .c_out(fc483));

	logic fs484, fc484;
	FA fa484 (.a(fc452), .b(fs475), .c_in(fs476), .s(fs484), .c_out(fc484));

	logic fs485, fc485;
	FA fa485 (.a(fs477), .b(fs478), .c_in(fc453), .s(fs485), .c_out(fc485));

	logic fs486, fc486;
	FA fa486 (.a(fs479), .b(fs480), .c_in(fs481), .s(fs486), .c_out(fc486));

	logic fs487, fc487;
	FA fa487 (.a(fc454), .b(fc455), .c_in(fc456), .s(fs487), .c_out(fc487));

	logic fs488, fc488;
	FA fa488 (.a(fs482), .b(fc457), .c_in(fs483), .s(fs488), .c_out(fc488));

	logic fs489, fc489;
	FA fa489 (.a(fs484), .b(fs485), .c_in(fc458), .s(fs489), .c_out(fc489));

	logic fs490, fc490;
	FA fa490 (.a(fs486), .b(fc459), .c_in(fc460), .s(fs490), .c_out(fc490));

	logic fs491, fc491;
	FA fa491 (.a(fs487), .b(fc461), .c_in(fs488), .s(fs491), .c_out(fc491));

	logic fs492, fc492;
	FA fa492 (.a(fs489), .b(fc462), .c_in(fs490), .s(fs492), .c_out(fc492));

	logic fs493, fc493;
	FA fa493 (.a(fc463), .b(fs491), .c_in(fs492), .s(fs493), .c_out(fc493));

	logic fs494, fc494;
	FA fa494 (.a(in_3_31), .b(in_4_30), .c_in(in_5_29), .s(fs494), .c_out(fc494));

	logic fs495, fc495;
	FA fa495 (.a(in_6_28), .b(in_7_27), .c_in(in_8_26), .s(fs495), .c_out(fc495));

	logic fs496, fc496;
	FA fa496 (.a(in_9_25), .b(in_10_24), .c_in(in_11_23), .s(fs496), .c_out(fc496));

	logic fs497, fc497;
	FA fa497 (.a(in_12_22), .b(in_13_21), .c_in(in_14_20), .s(fs497), .c_out(fc497));

	logic fs498, fc498;
	FA fa498 (.a(in_15_19), .b(in_16_18), .c_in(in_17_17), .s(fs498), .c_out(fc498));

	logic fs499, fc499;
	FA fa499 (.a(in_18_16), .b(in_19_15), .c_in(in_20_14), .s(fs499), .c_out(fc499));

	logic fs500, fc500;
	FA fa500 (.a(in_21_13), .b(in_22_12), .c_in(in_23_11), .s(fs500), .c_out(fc500));

	logic fs501, fc501;
	FA fa501 (.a(in_24_10), .b(in_25_9), .c_in(in_26_8), .s(fs501), .c_out(fc501));

	logic fs502, fc502;
	FA fa502 (.a(in_27_7), .b(in_28_6), .c_in(in_29_5), .s(fs502), .c_out(fc502));

	logic fs503, fc503;
	FA fa503 (.a(in_30_4), .b(in_31_3), .c_in(fc465), .s(fs503), .c_out(fc503));

	logic fs504, fc504;
	FA fa504 (.a(fc466), .b(fc467), .c_in(fc468), .s(fs504), .c_out(fc504));

	logic fs505, fc505;
	FA fa505 (.a(fc469), .b(fc470), .c_in(fc471), .s(fs505), .c_out(fc505));

	logic fs506, fc506;
	FA fa506 (.a(fc472), .b(fc473), .c_in(fc474), .s(fs506), .c_out(fc506));

	logic fs507, fc507;
	FA fa507 (.a(fs494), .b(fs495), .c_in(fs496), .s(fs507), .c_out(fc507));

	logic fs508, fc508;
	FA fa508 (.a(fs497), .b(fs498), .c_in(fs499), .s(fs508), .c_out(fc508));

	logic fs509, fc509;
	FA fa509 (.a(fs500), .b(fs501), .c_in(fs502), .s(fs509), .c_out(fc509));

	logic fs510, fc510;
	FA fa510 (.a(fc475), .b(fc476), .c_in(fc477), .s(fs510), .c_out(fc510));

	logic fs511, fc511;
	FA fa511 (.a(fc478), .b(fs503), .c_in(fc479), .s(fs511), .c_out(fc511));

	logic fs512, fc512;
	FA fa512 (.a(fc480), .b(fc481), .c_in(fs504), .s(fs512), .c_out(fc512));

	logic fs513, fc513;
	FA fa513 (.a(fs505), .b(fs506), .c_in(fc482), .s(fs513), .c_out(fc513));

	logic fs514, fc514;
	FA fa514 (.a(fs507), .b(fs508), .c_in(fs509), .s(fs514), .c_out(fc514));

	logic fs515, fc515;
	FA fa515 (.a(fc483), .b(fc484), .c_in(fc485), .s(fs515), .c_out(fc515));

	logic fs516, fc516;
	FA fa516 (.a(fs510), .b(fs511), .c_in(fc486), .s(fs516), .c_out(fc516));

	logic fs517, fc517;
	FA fa517 (.a(fs512), .b(fs513), .c_in(fc487), .s(fs517), .c_out(fc517));

	logic fs518, fc518;
	FA fa518 (.a(fs514), .b(fc488), .c_in(fc489), .s(fs518), .c_out(fc518));

	logic fs519, fc519;
	FA fa519 (.a(fs515), .b(fs516), .c_in(fs517), .s(fs519), .c_out(fc519));

	logic fs520, fc520;
	FA fa520 (.a(fc490), .b(fc491), .c_in(fs518), .s(fs520), .c_out(fc520));

	logic fs521, fc521;
	FA fa521 (.a(fs519), .b(fc492), .c_in(fs520), .s(fs521), .c_out(fc521));

	logic fs522, fc522;
	FA fa522 (.a(in_4_31), .b(in_5_30), .c_in(in_6_29), .s(fs522), .c_out(fc522));

	logic fs523, fc523;
	FA fa523 (.a(in_7_28), .b(in_8_27), .c_in(in_9_26), .s(fs523), .c_out(fc523));

	logic fs524, fc524;
	FA fa524 (.a(in_10_25), .b(in_11_24), .c_in(in_12_23), .s(fs524), .c_out(fc524));

	logic fs525, fc525;
	FA fa525 (.a(in_13_22), .b(in_14_21), .c_in(in_15_20), .s(fs525), .c_out(fc525));

	logic fs526, fc526;
	FA fa526 (.a(in_16_19), .b(in_17_18), .c_in(in_18_17), .s(fs526), .c_out(fc526));

	logic fs527, fc527;
	FA fa527 (.a(in_19_16), .b(in_20_15), .c_in(in_21_14), .s(fs527), .c_out(fc527));

	logic fs528, fc528;
	FA fa528 (.a(in_22_13), .b(in_23_12), .c_in(in_24_11), .s(fs528), .c_out(fc528));

	logic fs529, fc529;
	FA fa529 (.a(in_25_10), .b(in_26_9), .c_in(in_27_8), .s(fs529), .c_out(fc529));

	logic fs530, fc530;
	FA fa530 (.a(in_28_7), .b(in_29_6), .c_in(in_30_5), .s(fs530), .c_out(fc530));

	logic fs531, fc531;
	FA fa531 (.a(in_31_4), .b(fc494), .c_in(fc495), .s(fs531), .c_out(fc531));

	logic fs532, fc532;
	FA fa532 (.a(fc496), .b(fc497), .c_in(fc498), .s(fs532), .c_out(fc532));

	logic fs533, fc533;
	FA fa533 (.a(fc499), .b(fc500), .c_in(fc501), .s(fs533), .c_out(fc533));

	logic fs534, fc534;
	FA fa534 (.a(fc502), .b(fc503), .c_in(fs522), .s(fs534), .c_out(fc534));

	logic fs535, fc535;
	FA fa535 (.a(fs523), .b(fs524), .c_in(fs525), .s(fs535), .c_out(fc535));

	logic fs536, fc536;
	FA fa536 (.a(fs526), .b(fs527), .c_in(fs528), .s(fs536), .c_out(fc536));

	logic fs537, fc537;
	FA fa537 (.a(fs529), .b(fs530), .c_in(fc504), .s(fs537), .c_out(fc537));

	logic fs538, fc538;
	FA fa538 (.a(fc505), .b(fc506), .c_in(fc507), .s(fs538), .c_out(fc538));

	logic fs539, fc539;
	FA fa539 (.a(fc508), .b(fc509), .c_in(fs531), .s(fs539), .c_out(fc539));

	logic fs540, fc540;
	FA fa540 (.a(fs532), .b(fs533), .c_in(fc510), .s(fs540), .c_out(fc540));

	logic fs541, fc541;
	FA fa541 (.a(fc511), .b(fs534), .c_in(fs535), .s(fs541), .c_out(fc541));

	logic fs542, fc542;
	FA fa542 (.a(fs536), .b(fs537), .c_in(fc512), .s(fs542), .c_out(fc542));

	logic fs543, fc543;
	FA fa543 (.a(fc513), .b(fs538), .c_in(fc514), .s(fs543), .c_out(fc543));

	logic fs544, fc544;
	FA fa544 (.a(fs539), .b(fs540), .c_in(fc515), .s(fs544), .c_out(fc544));

	logic fs545, fc545;
	FA fa545 (.a(fc516), .b(fs541), .c_in(fs542), .s(fs545), .c_out(fc545));

	logic fs546, fc546;
	FA fa546 (.a(fc517), .b(fs543), .c_in(fs544), .s(fs546), .c_out(fc546));

	logic fs547, fc547;
	FA fa547 (.a(fc518), .b(fc519), .c_in(fs545), .s(fs547), .c_out(fc547));

	logic fs548, fc548;
	FA fa548 (.a(fs546), .b(fc520), .c_in(fs547), .s(fs548), .c_out(fc548));

	logic fs549, fc549;
	FA fa549 (.a(in_5_31), .b(in_6_30), .c_in(in_7_29), .s(fs549), .c_out(fc549));

	logic fs550, fc550;
	FA fa550 (.a(in_8_28), .b(in_9_27), .c_in(in_10_26), .s(fs550), .c_out(fc550));

	logic fs551, fc551;
	FA fa551 (.a(in_11_25), .b(in_12_24), .c_in(in_13_23), .s(fs551), .c_out(fc551));

	logic fs552, fc552;
	FA fa552 (.a(in_14_22), .b(in_15_21), .c_in(in_16_20), .s(fs552), .c_out(fc552));

	logic fs553, fc553;
	FA fa553 (.a(in_17_19), .b(in_18_18), .c_in(in_19_17), .s(fs553), .c_out(fc553));

	logic fs554, fc554;
	FA fa554 (.a(in_20_16), .b(in_21_15), .c_in(in_22_14), .s(fs554), .c_out(fc554));

	logic fs555, fc555;
	FA fa555 (.a(in_23_13), .b(in_24_12), .c_in(in_25_11), .s(fs555), .c_out(fc555));

	logic fs556, fc556;
	FA fa556 (.a(in_26_10), .b(in_27_9), .c_in(in_28_8), .s(fs556), .c_out(fc556));

	logic fs557, fc557;
	FA fa557 (.a(in_29_7), .b(in_30_6), .c_in(in_31_5), .s(fs557), .c_out(fc557));

	logic fs558, fc558;
	FA fa558 (.a(fc522), .b(fc523), .c_in(fc524), .s(fs558), .c_out(fc558));

	logic fs559, fc559;
	FA fa559 (.a(fc525), .b(fc526), .c_in(fc527), .s(fs559), .c_out(fc559));

	logic fs560, fc560;
	FA fa560 (.a(fc528), .b(fc529), .c_in(fc530), .s(fs560), .c_out(fc560));

	logic fs561, fc561;
	FA fa561 (.a(fs549), .b(fs550), .c_in(fs551), .s(fs561), .c_out(fc561));

	logic fs562, fc562;
	FA fa562 (.a(fs552), .b(fs553), .c_in(fs554), .s(fs562), .c_out(fc562));

	logic fs563, fc563;
	FA fa563 (.a(fs555), .b(fs556), .c_in(fs557), .s(fs563), .c_out(fc563));

	logic fs564, fc564;
	FA fa564 (.a(fc531), .b(fc532), .c_in(fc533), .s(fs564), .c_out(fc564));

	logic fs565, fc565;
	FA fa565 (.a(fc534), .b(fc535), .c_in(fc536), .s(fs565), .c_out(fc565));

	logic fs566, fc566;
	FA fa566 (.a(fc537), .b(fs558), .c_in(fs559), .s(fs566), .c_out(fc566));

	logic fs567, fc567;
	FA fa567 (.a(fs560), .b(fc538), .c_in(fs561), .s(fs567), .c_out(fc567));

	logic fs568, fc568;
	FA fa568 (.a(fs562), .b(fs563), .c_in(fc539), .s(fs568), .c_out(fc568));

	logic fs569, fc569;
	FA fa569 (.a(fc540), .b(fs564), .c_in(fc541), .s(fs569), .c_out(fc569));

	logic fs570, fc570;
	FA fa570 (.a(fc542), .b(fs565), .c_in(fs566), .s(fs570), .c_out(fc570));

	logic fs571, fc571;
	FA fa571 (.a(fc543), .b(fs567), .c_in(fs568), .s(fs571), .c_out(fc571));

	logic fs572, fc572;
	FA fa572 (.a(fc544), .b(fs569), .c_in(fc545), .s(fs572), .c_out(fc572));

	logic fs573, fc573;
	FA fa573 (.a(fs570), .b(fc546), .c_in(fs571), .s(fs573), .c_out(fc573));

	logic fs574, fc574;
	FA fa574 (.a(fs572), .b(fc547), .c_in(fs573), .s(fs574), .c_out(fc574));

	logic fs575, fc575;
	FA fa575 (.a(in_6_31), .b(in_7_30), .c_in(in_8_29), .s(fs575), .c_out(fc575));

	logic fs576, fc576;
	FA fa576 (.a(in_9_28), .b(in_10_27), .c_in(in_11_26), .s(fs576), .c_out(fc576));

	logic fs577, fc577;
	FA fa577 (.a(in_12_25), .b(in_13_24), .c_in(in_14_23), .s(fs577), .c_out(fc577));

	logic fs578, fc578;
	FA fa578 (.a(in_15_22), .b(in_16_21), .c_in(in_17_20), .s(fs578), .c_out(fc578));

	logic fs579, fc579;
	FA fa579 (.a(in_18_19), .b(in_19_18), .c_in(in_20_17), .s(fs579), .c_out(fc579));

	logic fs580, fc580;
	FA fa580 (.a(in_21_16), .b(in_22_15), .c_in(in_23_14), .s(fs580), .c_out(fc580));

	logic fs581, fc581;
	FA fa581 (.a(in_24_13), .b(in_25_12), .c_in(in_26_11), .s(fs581), .c_out(fc581));

	logic fs582, fc582;
	FA fa582 (.a(in_27_10), .b(in_28_9), .c_in(in_29_8), .s(fs582), .c_out(fc582));

	logic fs583, fc583;
	FA fa583 (.a(in_30_7), .b(in_31_6), .c_in(fc549), .s(fs583), .c_out(fc583));

	logic fs584, fc584;
	FA fa584 (.a(fc550), .b(fc551), .c_in(fc552), .s(fs584), .c_out(fc584));

	logic fs585, fc585;
	FA fa585 (.a(fc553), .b(fc554), .c_in(fc555), .s(fs585), .c_out(fc585));

	logic fs586, fc586;
	FA fa586 (.a(fc556), .b(fc557), .c_in(fs575), .s(fs586), .c_out(fc586));

	logic fs587, fc587;
	FA fa587 (.a(fs576), .b(fs577), .c_in(fs578), .s(fs587), .c_out(fc587));

	logic fs588, fc588;
	FA fa588 (.a(fs579), .b(fs580), .c_in(fs581), .s(fs588), .c_out(fc588));

	logic fs589, fc589;
	FA fa589 (.a(fs582), .b(fc558), .c_in(fc559), .s(fs589), .c_out(fc589));

	logic fs590, fc590;
	FA fa590 (.a(fc560), .b(fs583), .c_in(fc561), .s(fs590), .c_out(fc590));

	logic fs591, fc591;
	FA fa591 (.a(fc562), .b(fc563), .c_in(fs584), .s(fs591), .c_out(fc591));

	logic fs592, fc592;
	FA fa592 (.a(fs585), .b(fs586), .c_in(fc564), .s(fs592), .c_out(fc592));

	logic fs593, fc593;
	FA fa593 (.a(fs587), .b(fs588), .c_in(fc565), .s(fs593), .c_out(fc593));

	logic fs594, fc594;
	FA fa594 (.a(fc566), .b(fs589), .c_in(fs590), .s(fs594), .c_out(fc594));

	logic fs595, fc595;
	FA fa595 (.a(fc567), .b(fc568), .c_in(fs591), .s(fs595), .c_out(fc595));

	logic fs596, fc596;
	FA fa596 (.a(fs592), .b(fc569), .c_in(fs593), .s(fs596), .c_out(fc596));

	logic fs597, fc597;
	FA fa597 (.a(fc570), .b(fs594), .c_in(fc571), .s(fs597), .c_out(fc597));

	logic fs598, fc598;
	FA fa598 (.a(fs595), .b(fc572), .c_in(fs596), .s(fs598), .c_out(fc598));

	logic fs599, fc599;
	FA fa599 (.a(fs597), .b(fc573), .c_in(fs598), .s(fs599), .c_out(fc599));

	logic fs600, fc600;
	FA fa600 (.a(in_7_31), .b(in_8_30), .c_in(in_9_29), .s(fs600), .c_out(fc600));

	logic fs601, fc601;
	FA fa601 (.a(in_10_28), .b(in_11_27), .c_in(in_12_26), .s(fs601), .c_out(fc601));

	logic fs602, fc602;
	FA fa602 (.a(in_13_25), .b(in_14_24), .c_in(in_15_23), .s(fs602), .c_out(fc602));

	logic fs603, fc603;
	FA fa603 (.a(in_16_22), .b(in_17_21), .c_in(in_18_20), .s(fs603), .c_out(fc603));

	logic fs604, fc604;
	FA fa604 (.a(in_19_19), .b(in_20_18), .c_in(in_21_17), .s(fs604), .c_out(fc604));

	logic fs605, fc605;
	FA fa605 (.a(in_22_16), .b(in_23_15), .c_in(in_24_14), .s(fs605), .c_out(fc605));

	logic fs606, fc606;
	FA fa606 (.a(in_25_13), .b(in_26_12), .c_in(in_27_11), .s(fs606), .c_out(fc606));

	logic fs607, fc607;
	FA fa607 (.a(in_28_10), .b(in_29_9), .c_in(in_30_8), .s(fs607), .c_out(fc607));

	logic fs608, fc608;
	FA fa608 (.a(in_31_7), .b(fc575), .c_in(fc576), .s(fs608), .c_out(fc608));

	logic fs609, fc609;
	FA fa609 (.a(fc577), .b(fc578), .c_in(fc579), .s(fs609), .c_out(fc609));

	logic fs610, fc610;
	FA fa610 (.a(fc580), .b(fc581), .c_in(fc582), .s(fs610), .c_out(fc610));

	logic fs611, fc611;
	FA fa611 (.a(fc583), .b(fs600), .c_in(fs601), .s(fs611), .c_out(fc611));

	logic fs612, fc612;
	FA fa612 (.a(fs602), .b(fs603), .c_in(fs604), .s(fs612), .c_out(fc612));

	logic fs613, fc613;
	FA fa613 (.a(fs605), .b(fs606), .c_in(fs607), .s(fs613), .c_out(fc613));

	logic fs614, fc614;
	FA fa614 (.a(fc584), .b(fc585), .c_in(fc586), .s(fs614), .c_out(fc614));

	logic fs615, fc615;
	FA fa615 (.a(fc587), .b(fc588), .c_in(fs608), .s(fs615), .c_out(fc615));

	logic fs616, fc616;
	FA fa616 (.a(fs609), .b(fs610), .c_in(fc589), .s(fs616), .c_out(fc616));

	logic fs617, fc617;
	FA fa617 (.a(fc590), .b(fs611), .c_in(fs612), .s(fs617), .c_out(fc617));

	logic fs618, fc618;
	FA fa618 (.a(fs613), .b(fc591), .c_in(fc592), .s(fs618), .c_out(fc618));

	logic fs619, fc619;
	FA fa619 (.a(fs614), .b(fc593), .c_in(fs615), .s(fs619), .c_out(fc619));

	logic fs620, fc620;
	FA fa620 (.a(fs616), .b(fc594), .c_in(fs617), .s(fs620), .c_out(fc620));

	logic fs621, fc621;
	FA fa621 (.a(fc595), .b(fs618), .c_in(fc596), .s(fs621), .c_out(fc621));

	logic fs622, fc622;
	FA fa622 (.a(fs619), .b(fc597), .c_in(fs620), .s(fs622), .c_out(fc622));

	logic fs623, fc623;
	FA fa623 (.a(fs621), .b(fc598), .c_in(fs622), .s(fs623), .c_out(fc623));

	logic fs624, fc624;
	FA fa624 (.a(in_8_31), .b(in_9_30), .c_in(in_10_29), .s(fs624), .c_out(fc624));

	logic fs625, fc625;
	FA fa625 (.a(in_11_28), .b(in_12_27), .c_in(in_13_26), .s(fs625), .c_out(fc625));

	logic fs626, fc626;
	FA fa626 (.a(in_14_25), .b(in_15_24), .c_in(in_16_23), .s(fs626), .c_out(fc626));

	logic fs627, fc627;
	FA fa627 (.a(in_17_22), .b(in_18_21), .c_in(in_19_20), .s(fs627), .c_out(fc627));

	logic fs628, fc628;
	FA fa628 (.a(in_20_19), .b(in_21_18), .c_in(in_22_17), .s(fs628), .c_out(fc628));

	logic fs629, fc629;
	FA fa629 (.a(in_23_16), .b(in_24_15), .c_in(in_25_14), .s(fs629), .c_out(fc629));

	logic fs630, fc630;
	FA fa630 (.a(in_26_13), .b(in_27_12), .c_in(in_28_11), .s(fs630), .c_out(fc630));

	logic fs631, fc631;
	FA fa631 (.a(in_29_10), .b(in_30_9), .c_in(in_31_8), .s(fs631), .c_out(fc631));

	logic fs632, fc632;
	FA fa632 (.a(fc600), .b(fc601), .c_in(fc602), .s(fs632), .c_out(fc632));

	logic fs633, fc633;
	FA fa633 (.a(fc603), .b(fc604), .c_in(fc605), .s(fs633), .c_out(fc633));

	logic fs634, fc634;
	FA fa634 (.a(fc606), .b(fc607), .c_in(fs624), .s(fs634), .c_out(fc634));

	logic fs635, fc635;
	FA fa635 (.a(fs625), .b(fs626), .c_in(fs627), .s(fs635), .c_out(fc635));

	logic fs636, fc636;
	FA fa636 (.a(fs628), .b(fs629), .c_in(fs630), .s(fs636), .c_out(fc636));

	logic fs637, fc637;
	FA fa637 (.a(fs631), .b(fc608), .c_in(fc609), .s(fs637), .c_out(fc637));

	logic fs638, fc638;
	FA fa638 (.a(fc610), .b(fc611), .c_in(fc612), .s(fs638), .c_out(fc638));

	logic fs639, fc639;
	FA fa639 (.a(fc613), .b(fs632), .c_in(fs633), .s(fs639), .c_out(fc639));

	logic fs640, fc640;
	FA fa640 (.a(fs634), .b(fc614), .c_in(fs635), .s(fs640), .c_out(fc640));

	logic fs641, fc641;
	FA fa641 (.a(fs636), .b(fc615), .c_in(fc616), .s(fs641), .c_out(fc641));

	logic fs642, fc642;
	FA fa642 (.a(fs637), .b(fc617), .c_in(fs638), .s(fs642), .c_out(fc642));

	logic fs643, fc643;
	FA fa643 (.a(fs639), .b(fc618), .c_in(fs640), .s(fs643), .c_out(fc643));

	logic fs644, fc644;
	FA fa644 (.a(fc619), .b(fs641), .c_in(fc620), .s(fs644), .c_out(fc644));

	logic fs645, fc645;
	FA fa645 (.a(fs642), .b(fc621), .c_in(fs643), .s(fs645), .c_out(fc645));

	logic fs646, fc646;
	FA fa646 (.a(fs644), .b(fc622), .c_in(fs645), .s(fs646), .c_out(fc646));

	logic fs647, fc647;
	FA fa647 (.a(in_9_31), .b(in_10_30), .c_in(in_11_29), .s(fs647), .c_out(fc647));

	logic fs648, fc648;
	FA fa648 (.a(in_12_28), .b(in_13_27), .c_in(in_14_26), .s(fs648), .c_out(fc648));

	logic fs649, fc649;
	FA fa649 (.a(in_15_25), .b(in_16_24), .c_in(in_17_23), .s(fs649), .c_out(fc649));

	logic fs650, fc650;
	FA fa650 (.a(in_18_22), .b(in_19_21), .c_in(in_20_20), .s(fs650), .c_out(fc650));

	logic fs651, fc651;
	FA fa651 (.a(in_21_19), .b(in_22_18), .c_in(in_23_17), .s(fs651), .c_out(fc651));

	logic fs652, fc652;
	FA fa652 (.a(in_24_16), .b(in_25_15), .c_in(in_26_14), .s(fs652), .c_out(fc652));

	logic fs653, fc653;
	FA fa653 (.a(in_27_13), .b(in_28_12), .c_in(in_29_11), .s(fs653), .c_out(fc653));

	logic fs654, fc654;
	FA fa654 (.a(in_30_10), .b(in_31_9), .c_in(fc624), .s(fs654), .c_out(fc654));

	logic fs655, fc655;
	FA fa655 (.a(fc625), .b(fc626), .c_in(fc627), .s(fs655), .c_out(fc655));

	logic fs656, fc656;
	FA fa656 (.a(fc628), .b(fc629), .c_in(fc630), .s(fs656), .c_out(fc656));

	logic fs657, fc657;
	FA fa657 (.a(fc631), .b(fs647), .c_in(fs648), .s(fs657), .c_out(fc657));

	logic fs658, fc658;
	FA fa658 (.a(fs649), .b(fs650), .c_in(fs651), .s(fs658), .c_out(fc658));

	logic fs659, fc659;
	FA fa659 (.a(fs652), .b(fs653), .c_in(fc632), .s(fs659), .c_out(fc659));

	logic fs660, fc660;
	FA fa660 (.a(fc633), .b(fc634), .c_in(fs654), .s(fs660), .c_out(fc660));

	logic fs661, fc661;
	FA fa661 (.a(fc635), .b(fc636), .c_in(fs655), .s(fs661), .c_out(fc661));

	logic fs662, fc662;
	FA fa662 (.a(fs656), .b(fc637), .c_in(fs657), .s(fs662), .c_out(fc662));

	logic fs663, fc663;
	FA fa663 (.a(fs658), .b(fs659), .c_in(fc638), .s(fs663), .c_out(fc663));

	logic fs664, fc664;
	FA fa664 (.a(fc639), .b(fs660), .c_in(fc640), .s(fs664), .c_out(fc664));

	logic fs665, fc665;
	FA fa665 (.a(fs661), .b(fc641), .c_in(fs662), .s(fs665), .c_out(fc665));

	logic fs666, fc666;
	FA fa666 (.a(fs663), .b(fc642), .c_in(fs664), .s(fs666), .c_out(fc666));

	logic fs667, fc667;
	FA fa667 (.a(fc643), .b(fc644), .c_in(fs665), .s(fs667), .c_out(fc667));

	logic fs668, fc668;
	FA fa668 (.a(fs666), .b(fc645), .c_in(fs667), .s(fs668), .c_out(fc668));

	logic fs669, fc669;
	FA fa669 (.a(in_10_31), .b(in_11_30), .c_in(in_12_29), .s(fs669), .c_out(fc669));

	logic fs670, fc670;
	FA fa670 (.a(in_13_28), .b(in_14_27), .c_in(in_15_26), .s(fs670), .c_out(fc670));

	logic fs671, fc671;
	FA fa671 (.a(in_16_25), .b(in_17_24), .c_in(in_18_23), .s(fs671), .c_out(fc671));

	logic fs672, fc672;
	FA fa672 (.a(in_19_22), .b(in_20_21), .c_in(in_21_20), .s(fs672), .c_out(fc672));

	logic fs673, fc673;
	FA fa673 (.a(in_22_19), .b(in_23_18), .c_in(in_24_17), .s(fs673), .c_out(fc673));

	logic fs674, fc674;
	FA fa674 (.a(in_25_16), .b(in_26_15), .c_in(in_27_14), .s(fs674), .c_out(fc674));

	logic fs675, fc675;
	FA fa675 (.a(in_28_13), .b(in_29_12), .c_in(in_30_11), .s(fs675), .c_out(fc675));

	logic fs676, fc676;
	FA fa676 (.a(in_31_10), .b(fc647), .c_in(fc648), .s(fs676), .c_out(fc676));

	logic fs677, fc677;
	FA fa677 (.a(fc649), .b(fc650), .c_in(fc651), .s(fs677), .c_out(fc677));

	logic fs678, fc678;
	FA fa678 (.a(fc652), .b(fc653), .c_in(fc654), .s(fs678), .c_out(fc678));

	logic fs679, fc679;
	FA fa679 (.a(fs669), .b(fs670), .c_in(fs671), .s(fs679), .c_out(fc679));

	logic fs680, fc680;
	FA fa680 (.a(fs672), .b(fs673), .c_in(fs674), .s(fs680), .c_out(fc680));

	logic fs681, fc681;
	FA fa681 (.a(fs675), .b(fc655), .c_in(fc656), .s(fs681), .c_out(fc681));

	logic fs682, fc682;
	FA fa682 (.a(fc657), .b(fc658), .c_in(fc659), .s(fs682), .c_out(fc682));

	logic fs683, fc683;
	FA fa683 (.a(fs676), .b(fs677), .c_in(fs678), .s(fs683), .c_out(fc683));

	logic fs684, fc684;
	FA fa684 (.a(fc660), .b(fs679), .c_in(fs680), .s(fs684), .c_out(fc684));

	logic fs685, fc685;
	FA fa685 (.a(fc661), .b(fs681), .c_in(fc662), .s(fs685), .c_out(fc685));

	logic fs686, fc686;
	FA fa686 (.a(fc663), .b(fs682), .c_in(fs683), .s(fs686), .c_out(fc686));

	logic fs687, fc687;
	FA fa687 (.a(fc664), .b(fs684), .c_in(fs685), .s(fs687), .c_out(fc687));

	logic fs688, fc688;
	FA fa688 (.a(fc665), .b(fs686), .c_in(fc666), .s(fs688), .c_out(fc688));

	logic fs689, fc689;
	FA fa689 (.a(fs687), .b(fc667), .c_in(fs688), .s(fs689), .c_out(fc689));

	logic fs690, fc690;
	FA fa690 (.a(in_11_31), .b(in_12_30), .c_in(in_13_29), .s(fs690), .c_out(fc690));

	logic fs691, fc691;
	FA fa691 (.a(in_14_28), .b(in_15_27), .c_in(in_16_26), .s(fs691), .c_out(fc691));

	logic fs692, fc692;
	FA fa692 (.a(in_17_25), .b(in_18_24), .c_in(in_19_23), .s(fs692), .c_out(fc692));

	logic fs693, fc693;
	FA fa693 (.a(in_20_22), .b(in_21_21), .c_in(in_22_20), .s(fs693), .c_out(fc693));

	logic fs694, fc694;
	FA fa694 (.a(in_23_19), .b(in_24_18), .c_in(in_25_17), .s(fs694), .c_out(fc694));

	logic fs695, fc695;
	FA fa695 (.a(in_26_16), .b(in_27_15), .c_in(in_28_14), .s(fs695), .c_out(fc695));

	logic fs696, fc696;
	FA fa696 (.a(in_29_13), .b(in_30_12), .c_in(in_31_11), .s(fs696), .c_out(fc696));

	logic fs697, fc697;
	FA fa697 (.a(fc669), .b(fc670), .c_in(fc671), .s(fs697), .c_out(fc697));

	logic fs698, fc698;
	FA fa698 (.a(fc672), .b(fc673), .c_in(fc674), .s(fs698), .c_out(fc698));

	logic fs699, fc699;
	FA fa699 (.a(fc675), .b(fs690), .c_in(fs691), .s(fs699), .c_out(fc699));

	logic fs700, fc700;
	FA fa700 (.a(fs692), .b(fs693), .c_in(fs694), .s(fs700), .c_out(fc700));

	logic fs701, fc701;
	FA fa701 (.a(fs695), .b(fs696), .c_in(fc676), .s(fs701), .c_out(fc701));

	logic fs702, fc702;
	FA fa702 (.a(fc677), .b(fc678), .c_in(fc679), .s(fs702), .c_out(fc702));

	logic fs703, fc703;
	FA fa703 (.a(fc680), .b(fs697), .c_in(fs698), .s(fs703), .c_out(fc703));

	logic fs704, fc704;
	FA fa704 (.a(fc681), .b(fs699), .c_in(fs700), .s(fs704), .c_out(fc704));

	logic fs705, fc705;
	FA fa705 (.a(fs701), .b(fc682), .c_in(fc683), .s(fs705), .c_out(fc705));

	logic fs706, fc706;
	FA fa706 (.a(fs702), .b(fc684), .c_in(fs703), .s(fs706), .c_out(fc706));

	logic fs707, fc707;
	FA fa707 (.a(fc685), .b(fs704), .c_in(fc686), .s(fs707), .c_out(fc707));

	logic fs708, fc708;
	FA fa708 (.a(fs705), .b(fc687), .c_in(fs706), .s(fs708), .c_out(fc708));

	logic fs709, fc709;
	FA fa709 (.a(fs707), .b(fc688), .c_in(fs708), .s(fs709), .c_out(fc709));

	logic fs710, fc710;
	FA fa710 (.a(in_12_31), .b(in_13_30), .c_in(in_14_29), .s(fs710), .c_out(fc710));

	logic fs711, fc711;
	FA fa711 (.a(in_15_28), .b(in_16_27), .c_in(in_17_26), .s(fs711), .c_out(fc711));

	logic fs712, fc712;
	FA fa712 (.a(in_18_25), .b(in_19_24), .c_in(in_20_23), .s(fs712), .c_out(fc712));

	logic fs713, fc713;
	FA fa713 (.a(in_21_22), .b(in_22_21), .c_in(in_23_20), .s(fs713), .c_out(fc713));

	logic fs714, fc714;
	FA fa714 (.a(in_24_19), .b(in_25_18), .c_in(in_26_17), .s(fs714), .c_out(fc714));

	logic fs715, fc715;
	FA fa715 (.a(in_27_16), .b(in_28_15), .c_in(in_29_14), .s(fs715), .c_out(fc715));

	logic fs716, fc716;
	FA fa716 (.a(in_30_13), .b(in_31_12), .c_in(fc690), .s(fs716), .c_out(fc716));

	logic fs717, fc717;
	FA fa717 (.a(fc691), .b(fc692), .c_in(fc693), .s(fs717), .c_out(fc717));

	logic fs718, fc718;
	FA fa718 (.a(fc694), .b(fc695), .c_in(fc696), .s(fs718), .c_out(fc718));

	logic fs719, fc719;
	FA fa719 (.a(fs710), .b(fs711), .c_in(fs712), .s(fs719), .c_out(fc719));

	logic fs720, fc720;
	FA fa720 (.a(fs713), .b(fs714), .c_in(fs715), .s(fs720), .c_out(fc720));

	logic fs721, fc721;
	FA fa721 (.a(fc697), .b(fc698), .c_in(fs716), .s(fs721), .c_out(fc721));

	logic fs722, fc722;
	FA fa722 (.a(fc699), .b(fc700), .c_in(fc701), .s(fs722), .c_out(fc722));

	logic fs723, fc723;
	FA fa723 (.a(fs717), .b(fs718), .c_in(fc702), .s(fs723), .c_out(fc723));

	logic fs724, fc724;
	FA fa724 (.a(fs719), .b(fs720), .c_in(fc703), .s(fs724), .c_out(fc724));

	logic fs725, fc725;
	FA fa725 (.a(fs721), .b(fc704), .c_in(fs722), .s(fs725), .c_out(fc725));

	logic fs726, fc726;
	FA fa726 (.a(fs723), .b(fc705), .c_in(fs724), .s(fs726), .c_out(fc726));

	logic fs727, fc727;
	FA fa727 (.a(fc706), .b(fc707), .c_in(fs725), .s(fs727), .c_out(fc727));

	logic fs728, fc728;
	FA fa728 (.a(fs726), .b(fc708), .c_in(fs727), .s(fs728), .c_out(fc728));

	logic fs729, fc729;
	FA fa729 (.a(in_13_31), .b(in_14_30), .c_in(in_15_29), .s(fs729), .c_out(fc729));

	logic fs730, fc730;
	FA fa730 (.a(in_16_28), .b(in_17_27), .c_in(in_18_26), .s(fs730), .c_out(fc730));

	logic fs731, fc731;
	FA fa731 (.a(in_19_25), .b(in_20_24), .c_in(in_21_23), .s(fs731), .c_out(fc731));

	logic fs732, fc732;
	FA fa732 (.a(in_22_22), .b(in_23_21), .c_in(in_24_20), .s(fs732), .c_out(fc732));

	logic fs733, fc733;
	FA fa733 (.a(in_25_19), .b(in_26_18), .c_in(in_27_17), .s(fs733), .c_out(fc733));

	logic fs734, fc734;
	FA fa734 (.a(in_28_16), .b(in_29_15), .c_in(in_30_14), .s(fs734), .c_out(fc734));

	logic fs735, fc735;
	FA fa735 (.a(in_31_13), .b(fc710), .c_in(fc711), .s(fs735), .c_out(fc735));

	logic fs736, fc736;
	FA fa736 (.a(fc712), .b(fc713), .c_in(fc714), .s(fs736), .c_out(fc736));

	logic fs737, fc737;
	FA fa737 (.a(fc715), .b(fc716), .c_in(fs729), .s(fs737), .c_out(fc737));

	logic fs738, fc738;
	FA fa738 (.a(fs730), .b(fs731), .c_in(fs732), .s(fs738), .c_out(fc738));

	logic fs739, fc739;
	FA fa739 (.a(fs733), .b(fs734), .c_in(fc717), .s(fs739), .c_out(fc739));

	logic fs740, fc740;
	FA fa740 (.a(fc718), .b(fc719), .c_in(fc720), .s(fs740), .c_out(fc740));

	logic fs741, fc741;
	FA fa741 (.a(fs735), .b(fs736), .c_in(fc721), .s(fs741), .c_out(fc741));

	logic fs742, fc742;
	FA fa742 (.a(fs737), .b(fs738), .c_in(fs739), .s(fs742), .c_out(fc742));

	logic fs743, fc743;
	FA fa743 (.a(fc722), .b(fc723), .c_in(fc724), .s(fs743), .c_out(fc743));

	logic fs744, fc744;
	FA fa744 (.a(fs740), .b(fs741), .c_in(fs742), .s(fs744), .c_out(fc744));

	logic fs745, fc745;
	FA fa745 (.a(fc725), .b(fs743), .c_in(fc726), .s(fs745), .c_out(fc745));

	logic fs746, fc746;
	FA fa746 (.a(fs744), .b(fc727), .c_in(fs745), .s(fs746), .c_out(fc746));

	logic fs747, fc747;
	FA fa747 (.a(in_14_31), .b(in_15_30), .c_in(in_16_29), .s(fs747), .c_out(fc747));

	logic fs748, fc748;
	FA fa748 (.a(in_17_28), .b(in_18_27), .c_in(in_19_26), .s(fs748), .c_out(fc748));

	logic fs749, fc749;
	FA fa749 (.a(in_20_25), .b(in_21_24), .c_in(in_22_23), .s(fs749), .c_out(fc749));

	logic fs750, fc750;
	FA fa750 (.a(in_23_22), .b(in_24_21), .c_in(in_25_20), .s(fs750), .c_out(fc750));

	logic fs751, fc751;
	FA fa751 (.a(in_26_19), .b(in_27_18), .c_in(in_28_17), .s(fs751), .c_out(fc751));

	logic fs752, fc752;
	FA fa752 (.a(in_29_16), .b(in_30_15), .c_in(in_31_14), .s(fs752), .c_out(fc752));

	logic fs753, fc753;
	FA fa753 (.a(fc729), .b(fc730), .c_in(fc731), .s(fs753), .c_out(fc753));

	logic fs754, fc754;
	FA fa754 (.a(fc732), .b(fc733), .c_in(fc734), .s(fs754), .c_out(fc754));

	logic fs755, fc755;
	FA fa755 (.a(fs747), .b(fs748), .c_in(fs749), .s(fs755), .c_out(fc755));

	logic fs756, fc756;
	FA fa756 (.a(fs750), .b(fs751), .c_in(fs752), .s(fs756), .c_out(fc756));

	logic fs757, fc757;
	FA fa757 (.a(fc735), .b(fc736), .c_in(fc737), .s(fs757), .c_out(fc757));

	logic fs758, fc758;
	FA fa758 (.a(fc738), .b(fc739), .c_in(fs753), .s(fs758), .c_out(fc758));

	logic fs759, fc759;
	FA fa759 (.a(fs754), .b(fs755), .c_in(fs756), .s(fs759), .c_out(fc759));

	logic fs760, fc760;
	FA fa760 (.a(fc740), .b(fc741), .c_in(fs757), .s(fs760), .c_out(fc760));

	logic fs761, fc761;
	FA fa761 (.a(fc742), .b(fs758), .c_in(fc743), .s(fs761), .c_out(fc761));

	logic fs762, fc762;
	FA fa762 (.a(fs759), .b(fc744), .c_in(fs760), .s(fs762), .c_out(fc762));

	logic fs763, fc763;
	FA fa763 (.a(fs761), .b(fc745), .c_in(fs762), .s(fs763), .c_out(fc763));

	logic fs764, fc764;
	FA fa764 (.a(in_15_31), .b(in_16_30), .c_in(in_17_29), .s(fs764), .c_out(fc764));

	logic fs765, fc765;
	FA fa765 (.a(in_18_28), .b(in_19_27), .c_in(in_20_26), .s(fs765), .c_out(fc765));

	logic fs766, fc766;
	FA fa766 (.a(in_21_25), .b(in_22_24), .c_in(in_23_23), .s(fs766), .c_out(fc766));

	logic fs767, fc767;
	FA fa767 (.a(in_24_22), .b(in_25_21), .c_in(in_26_20), .s(fs767), .c_out(fc767));

	logic fs768, fc768;
	FA fa768 (.a(in_27_19), .b(in_28_18), .c_in(in_29_17), .s(fs768), .c_out(fc768));

	logic fs769, fc769;
	FA fa769 (.a(in_30_16), .b(in_31_15), .c_in(fc747), .s(fs769), .c_out(fc769));

	logic fs770, fc770;
	FA fa770 (.a(fc748), .b(fc749), .c_in(fc750), .s(fs770), .c_out(fc770));

	logic fs771, fc771;
	FA fa771 (.a(fc751), .b(fc752), .c_in(fs764), .s(fs771), .c_out(fc771));

	logic fs772, fc772;
	FA fa772 (.a(fs765), .b(fs766), .c_in(fs767), .s(fs772), .c_out(fc772));

	logic fs773, fc773;
	FA fa773 (.a(fs768), .b(fc753), .c_in(fc754), .s(fs773), .c_out(fc773));

	logic fs774, fc774;
	FA fa774 (.a(fs769), .b(fc755), .c_in(fc756), .s(fs774), .c_out(fc774));

	logic fs775, fc775;
	FA fa775 (.a(fs770), .b(fs771), .c_in(fc757), .s(fs775), .c_out(fc775));

	logic fs776, fc776;
	FA fa776 (.a(fs772), .b(fc758), .c_in(fs773), .s(fs776), .c_out(fc776));

	logic fs777, fc777;
	FA fa777 (.a(fc759), .b(fs774), .c_in(fs775), .s(fs777), .c_out(fc777));

	logic fs778, fc778;
	FA fa778 (.a(fc760), .b(fc761), .c_in(fs776), .s(fs778), .c_out(fc778));

	logic fs779, fc779;
	FA fa779 (.a(fs777), .b(fc762), .c_in(fs778), .s(fs779), .c_out(fc779));

	logic fs780, fc780;
	FA fa780 (.a(in_16_31), .b(in_17_30), .c_in(in_18_29), .s(fs780), .c_out(fc780));

	logic fs781, fc781;
	FA fa781 (.a(in_19_28), .b(in_20_27), .c_in(in_21_26), .s(fs781), .c_out(fc781));

	logic fs782, fc782;
	FA fa782 (.a(in_22_25), .b(in_23_24), .c_in(in_24_23), .s(fs782), .c_out(fc782));

	logic fs783, fc783;
	FA fa783 (.a(in_25_22), .b(in_26_21), .c_in(in_27_20), .s(fs783), .c_out(fc783));

	logic fs784, fc784;
	FA fa784 (.a(in_28_19), .b(in_29_18), .c_in(in_30_17), .s(fs784), .c_out(fc784));

	logic fs785, fc785;
	FA fa785 (.a(in_31_16), .b(fc764), .c_in(fc765), .s(fs785), .c_out(fc785));

	logic fs786, fc786;
	FA fa786 (.a(fc766), .b(fc767), .c_in(fc768), .s(fs786), .c_out(fc786));

	logic fs787, fc787;
	FA fa787 (.a(fc769), .b(fs780), .c_in(fs781), .s(fs787), .c_out(fc787));

	logic fs788, fc788;
	FA fa788 (.a(fs782), .b(fs783), .c_in(fs784), .s(fs788), .c_out(fc788));

	logic fs789, fc789;
	FA fa789 (.a(fc770), .b(fc771), .c_in(fc772), .s(fs789), .c_out(fc789));

	logic fs790, fc790;
	FA fa790 (.a(fs785), .b(fs786), .c_in(fc773), .s(fs790), .c_out(fc790));

	logic fs791, fc791;
	FA fa791 (.a(fs787), .b(fs788), .c_in(fc774), .s(fs791), .c_out(fc791));

	logic fs792, fc792;
	FA fa792 (.a(fc775), .b(fs789), .c_in(fs790), .s(fs792), .c_out(fc792));

	logic fs793, fc793;
	FA fa793 (.a(fc776), .b(fs791), .c_in(fc777), .s(fs793), .c_out(fc793));

	logic fs794, fc794;
	FA fa794 (.a(fs792), .b(fc778), .c_in(fs793), .s(fs794), .c_out(fc794));

	logic fs795, fc795;
	FA fa795 (.a(in_17_31), .b(in_18_30), .c_in(in_19_29), .s(fs795), .c_out(fc795));

	logic fs796, fc796;
	FA fa796 (.a(in_20_28), .b(in_21_27), .c_in(in_22_26), .s(fs796), .c_out(fc796));

	logic fs797, fc797;
	FA fa797 (.a(in_23_25), .b(in_24_24), .c_in(in_25_23), .s(fs797), .c_out(fc797));

	logic fs798, fc798;
	FA fa798 (.a(in_26_22), .b(in_27_21), .c_in(in_28_20), .s(fs798), .c_out(fc798));

	logic fs799, fc799;
	FA fa799 (.a(in_29_19), .b(in_30_18), .c_in(in_31_17), .s(fs799), .c_out(fc799));

	logic fs800, fc800;
	FA fa800 (.a(fc780), .b(fc781), .c_in(fc782), .s(fs800), .c_out(fc800));

	logic fs801, fc801;
	FA fa801 (.a(fc783), .b(fc784), .c_in(fs795), .s(fs801), .c_out(fc801));

	logic fs802, fc802;
	FA fa802 (.a(fs796), .b(fs797), .c_in(fs798), .s(fs802), .c_out(fc802));

	logic fs803, fc803;
	FA fa803 (.a(fs799), .b(fc785), .c_in(fc786), .s(fs803), .c_out(fc803));

	logic fs804, fc804;
	FA fa804 (.a(fc787), .b(fc788), .c_in(fs800), .s(fs804), .c_out(fc804));

	logic fs805, fc805;
	FA fa805 (.a(fs801), .b(fc789), .c_in(fs802), .s(fs805), .c_out(fc805));

	logic fs806, fc806;
	FA fa806 (.a(fc790), .b(fs803), .c_in(fc791), .s(fs806), .c_out(fc806));

	logic fs807, fc807;
	FA fa807 (.a(fs804), .b(fc792), .c_in(fs805), .s(fs807), .c_out(fc807));

	logic fs808, fc808;
	FA fa808 (.a(fs806), .b(fc793), .c_in(fs807), .s(fs808), .c_out(fc808));

	logic fs809, fc809;
	FA fa809 (.a(in_18_31), .b(in_19_30), .c_in(in_20_29), .s(fs809), .c_out(fc809));

	logic fs810, fc810;
	FA fa810 (.a(in_21_28), .b(in_22_27), .c_in(in_23_26), .s(fs810), .c_out(fc810));

	logic fs811, fc811;
	FA fa811 (.a(in_24_25), .b(in_25_24), .c_in(in_26_23), .s(fs811), .c_out(fc811));

	logic fs812, fc812;
	FA fa812 (.a(in_27_22), .b(in_28_21), .c_in(in_29_20), .s(fs812), .c_out(fc812));

	logic fs813, fc813;
	FA fa813 (.a(in_30_19), .b(in_31_18), .c_in(fc795), .s(fs813), .c_out(fc813));

	logic fs814, fc814;
	FA fa814 (.a(fc796), .b(fc797), .c_in(fc798), .s(fs814), .c_out(fc814));

	logic fs815, fc815;
	FA fa815 (.a(fc799), .b(fs809), .c_in(fs810), .s(fs815), .c_out(fc815));

	logic fs816, fc816;
	FA fa816 (.a(fs811), .b(fs812), .c_in(fc800), .s(fs816), .c_out(fc816));

	logic fs817, fc817;
	FA fa817 (.a(fc801), .b(fs813), .c_in(fc802), .s(fs817), .c_out(fc817));

	logic fs818, fc818;
	FA fa818 (.a(fs814), .b(fc803), .c_in(fs815), .s(fs818), .c_out(fc818));

	logic fs819, fc819;
	FA fa819 (.a(fs816), .b(fc804), .c_in(fs817), .s(fs819), .c_out(fc819));

	logic fs820, fc820;
	FA fa820 (.a(fc805), .b(fc806), .c_in(fs818), .s(fs820), .c_out(fc820));

	logic fs821, fc821;
	FA fa821 (.a(fs819), .b(fc807), .c_in(fs820), .s(fs821), .c_out(fc821));

	logic fs822, fc822;
	FA fa822 (.a(in_19_31), .b(in_20_30), .c_in(in_21_29), .s(fs822), .c_out(fc822));

	logic fs823, fc823;
	FA fa823 (.a(in_22_28), .b(in_23_27), .c_in(in_24_26), .s(fs823), .c_out(fc823));

	logic fs824, fc824;
	FA fa824 (.a(in_25_25), .b(in_26_24), .c_in(in_27_23), .s(fs824), .c_out(fc824));

	logic fs825, fc825;
	FA fa825 (.a(in_28_22), .b(in_29_21), .c_in(in_30_20), .s(fs825), .c_out(fc825));

	logic fs826, fc826;
	FA fa826 (.a(in_31_19), .b(fc809), .c_in(fc810), .s(fs826), .c_out(fc826));

	logic fs827, fc827;
	FA fa827 (.a(fc811), .b(fc812), .c_in(fc813), .s(fs827), .c_out(fc827));

	logic fs828, fc828;
	FA fa828 (.a(fs822), .b(fs823), .c_in(fs824), .s(fs828), .c_out(fc828));

	logic fs829, fc829;
	FA fa829 (.a(fs825), .b(fc814), .c_in(fc815), .s(fs829), .c_out(fc829));

	logic fs830, fc830;
	FA fa830 (.a(fc816), .b(fs826), .c_in(fs827), .s(fs830), .c_out(fc830));

	logic fs831, fc831;
	FA fa831 (.a(fc817), .b(fs828), .c_in(fs829), .s(fs831), .c_out(fc831));

	logic fs832, fc832;
	FA fa832 (.a(fc818), .b(fs830), .c_in(fc819), .s(fs832), .c_out(fc832));

	logic fs833, fc833;
	FA fa833 (.a(fs831), .b(fc820), .c_in(fs832), .s(fs833), .c_out(fc833));

	logic fs834, fc834;
	FA fa834 (.a(in_20_31), .b(in_21_30), .c_in(in_22_29), .s(fs834), .c_out(fc834));

	logic fs835, fc835;
	FA fa835 (.a(in_23_28), .b(in_24_27), .c_in(in_25_26), .s(fs835), .c_out(fc835));

	logic fs836, fc836;
	FA fa836 (.a(in_26_25), .b(in_27_24), .c_in(in_28_23), .s(fs836), .c_out(fc836));

	logic fs837, fc837;
	FA fa837 (.a(in_29_22), .b(in_30_21), .c_in(in_31_20), .s(fs837), .c_out(fc837));

	logic fs838, fc838;
	FA fa838 (.a(fc822), .b(fc823), .c_in(fc824), .s(fs838), .c_out(fc838));

	logic fs839, fc839;
	FA fa839 (.a(fc825), .b(fs834), .c_in(fs835), .s(fs839), .c_out(fc839));

	logic fs840, fc840;
	FA fa840 (.a(fs836), .b(fs837), .c_in(fc826), .s(fs840), .c_out(fc840));

	logic fs841, fc841;
	FA fa841 (.a(fc827), .b(fc828), .c_in(fs838), .s(fs841), .c_out(fc841));

	logic fs842, fc842;
	FA fa842 (.a(fc829), .b(fs839), .c_in(fs840), .s(fs842), .c_out(fc842));

	logic fs843, fc843;
	FA fa843 (.a(fc830), .b(fc831), .c_in(fs841), .s(fs843), .c_out(fc843));

	logic fs844, fc844;
	FA fa844 (.a(fs842), .b(fc832), .c_in(fs843), .s(fs844), .c_out(fc844));

	logic fs845, fc845;
	FA fa845 (.a(in_21_31), .b(in_22_30), .c_in(in_23_29), .s(fs845), .c_out(fc845));

	logic fs846, fc846;
	FA fa846 (.a(in_24_28), .b(in_25_27), .c_in(in_26_26), .s(fs846), .c_out(fc846));

	logic fs847, fc847;
	FA fa847 (.a(in_27_25), .b(in_28_24), .c_in(in_29_23), .s(fs847), .c_out(fc847));

	logic fs848, fc848;
	FA fa848 (.a(in_30_22), .b(in_31_21), .c_in(fc834), .s(fs848), .c_out(fc848));

	logic fs849, fc849;
	FA fa849 (.a(fc835), .b(fc836), .c_in(fc837), .s(fs849), .c_out(fc849));

	logic fs850, fc850;
	FA fa850 (.a(fs845), .b(fs846), .c_in(fs847), .s(fs850), .c_out(fc850));

	logic fs851, fc851;
	FA fa851 (.a(fc838), .b(fs848), .c_in(fc839), .s(fs851), .c_out(fc851));

	logic fs852, fc852;
	FA fa852 (.a(fc840), .b(fs849), .c_in(fs850), .s(fs852), .c_out(fc852));

	logic fs853, fc853;
	FA fa853 (.a(fc841), .b(fs851), .c_in(fc842), .s(fs853), .c_out(fc853));

	logic fs854, fc854;
	FA fa854 (.a(fs852), .b(fc843), .c_in(fs853), .s(fs854), .c_out(fc854));

	logic fs855, fc855;
	FA fa855 (.a(in_22_31), .b(in_23_30), .c_in(in_24_29), .s(fs855), .c_out(fc855));

	logic fs856, fc856;
	FA fa856 (.a(in_25_28), .b(in_26_27), .c_in(in_27_26), .s(fs856), .c_out(fc856));

	logic fs857, fc857;
	FA fa857 (.a(in_28_25), .b(in_29_24), .c_in(in_30_23), .s(fs857), .c_out(fc857));

	logic fs858, fc858;
	FA fa858 (.a(in_31_22), .b(fc845), .c_in(fc846), .s(fs858), .c_out(fc858));

	logic fs859, fc859;
	FA fa859 (.a(fc847), .b(fc848), .c_in(fs855), .s(fs859), .c_out(fc859));

	logic fs860, fc860;
	FA fa860 (.a(fs856), .b(fs857), .c_in(fc849), .s(fs860), .c_out(fc860));

	logic fs861, fc861;
	FA fa861 (.a(fc850), .b(fs858), .c_in(fc851), .s(fs861), .c_out(fc861));

	logic fs862, fc862;
	FA fa862 (.a(fs859), .b(fs860), .c_in(fc852), .s(fs862), .c_out(fc862));

	logic fs863, fc863;
	FA fa863 (.a(fs861), .b(fc853), .c_in(fs862), .s(fs863), .c_out(fc863));

	logic fs864, fc864;
	FA fa864 (.a(in_23_31), .b(in_24_30), .c_in(in_25_29), .s(fs864), .c_out(fc864));

	logic fs865, fc865;
	FA fa865 (.a(in_26_28), .b(in_27_27), .c_in(in_28_26), .s(fs865), .c_out(fc865));

	logic fs866, fc866;
	FA fa866 (.a(in_29_25), .b(in_30_24), .c_in(in_31_23), .s(fs866), .c_out(fc866));

	logic fs867, fc867;
	FA fa867 (.a(fc855), .b(fc856), .c_in(fc857), .s(fs867), .c_out(fc867));

	logic fs868, fc868;
	FA fa868 (.a(fs864), .b(fs865), .c_in(fs866), .s(fs868), .c_out(fc868));

	logic fs869, fc869;
	FA fa869 (.a(fc858), .b(fc859), .c_in(fc860), .s(fs869), .c_out(fc869));

	logic fs870, fc870;
	FA fa870 (.a(fs867), .b(fs868), .c_in(fc861), .s(fs870), .c_out(fc870));

	logic fs871, fc871;
	FA fa871 (.a(fc862), .b(fs869), .c_in(fs870), .s(fs871), .c_out(fc871));

	logic fs872, fc872;
	FA fa872 (.a(in_24_31), .b(in_25_30), .c_in(in_26_29), .s(fs872), .c_out(fc872));

	logic fs873, fc873;
	FA fa873 (.a(in_27_28), .b(in_28_27), .c_in(in_29_26), .s(fs873), .c_out(fc873));

	logic fs874, fc874;
	FA fa874 (.a(in_30_25), .b(in_31_24), .c_in(fc864), .s(fs874), .c_out(fc874));

	logic fs875, fc875;
	FA fa875 (.a(fc865), .b(fc866), .c_in(fs872), .s(fs875), .c_out(fc875));

	logic fs876, fc876;
	FA fa876 (.a(fs873), .b(fc867), .c_in(fs874), .s(fs876), .c_out(fc876));

	logic fs877, fc877;
	FA fa877 (.a(fc868), .b(fs875), .c_in(fc869), .s(fs877), .c_out(fc877));

	logic fs878, fc878;
	FA fa878 (.a(fs876), .b(fc870), .c_in(fs877), .s(fs878), .c_out(fc878));

	logic fs879, fc879;
	FA fa879 (.a(in_25_31), .b(in_26_30), .c_in(in_27_29), .s(fs879), .c_out(fc879));

	logic fs880, fc880;
	FA fa880 (.a(in_28_28), .b(in_29_27), .c_in(in_30_26), .s(fs880), .c_out(fc880));

	logic fs881, fc881;
	FA fa881 (.a(in_31_25), .b(fc872), .c_in(fc873), .s(fs881), .c_out(fc881));

	logic fs882, fc882;
	FA fa882 (.a(fc874), .b(fs879), .c_in(fs880), .s(fs882), .c_out(fc882));

	logic fs883, fc883;
	FA fa883 (.a(fc875), .b(fs881), .c_in(fc876), .s(fs883), .c_out(fc883));

	logic fs884, fc884;
	FA fa884 (.a(fs882), .b(fc877), .c_in(fs883), .s(fs884), .c_out(fc884));

	logic fs885, fc885;
	FA fa885 (.a(in_26_31), .b(in_27_30), .c_in(in_28_29), .s(fs885), .c_out(fc885));

	logic fs886, fc886;
	FA fa886 (.a(in_29_28), .b(in_30_27), .c_in(in_31_26), .s(fs886), .c_out(fc886));

	logic fs887, fc887;
	FA fa887 (.a(fc879), .b(fc880), .c_in(fs885), .s(fs887), .c_out(fc887));

	logic fs888, fc888;
	FA fa888 (.a(fs886), .b(fc881), .c_in(fc882), .s(fs888), .c_out(fc888));

	logic fs889, fc889;
	FA fa889 (.a(fs887), .b(fc883), .c_in(fs888), .s(fs889), .c_out(fc889));

	logic fs890, fc890;
	FA fa890 (.a(in_27_31), .b(in_28_30), .c_in(in_29_29), .s(fs890), .c_out(fc890));

	logic fs891, fc891;
	FA fa891 (.a(in_30_28), .b(in_31_27), .c_in(fc885), .s(fs891), .c_out(fc891));

	logic fs892, fc892;
	FA fa892 (.a(fc886), .b(fs890), .c_in(fc887), .s(fs892), .c_out(fc892));

	logic fs893, fc893;
	FA fa893 (.a(fs891), .b(fc888), .c_in(fs892), .s(fs893), .c_out(fc893));

	logic fs894, fc894;
	FA fa894 (.a(in_28_31), .b(in_29_30), .c_in(in_30_29), .s(fs894), .c_out(fc894));

	logic fs895, fc895;
	FA fa895 (.a(in_31_28), .b(fc890), .c_in(fc891), .s(fs895), .c_out(fc895));

	logic fs896, fc896;
	FA fa896 (.a(fs894), .b(fc892), .c_in(fs895), .s(fs896), .c_out(fc896));

	logic fs897, fc897;
	FA fa897 (.a(in_29_31), .b(in_30_30), .c_in(in_31_29), .s(fs897), .c_out(fc897));

	logic fs898, fc898;
	FA fa898 (.a(fc894), .b(fc895), .c_in(fs897), .s(fs898), .c_out(fc898));

	logic fs899, fc899;
	FA fa899 (.a(in_30_31), .b(in_31_30), .c_in(fc897), .s(fs899), .c_out(fc899));

	logic[62:0] cpa0, cpa1;

	assign cpa0 = {in_31_31, fc898, fc896, fc893, fc889, fc884, fc878, fc871, fc863, fc854, fc844, fc833, fc821, fc808, fc794, fc779, fc763, fc746, fc728, fc709, fc689, fc668, fc646, fc623, fc599, fc574, fc548, fc521, fc493, fc464, fc435, fc406, fc378, fc351, fc325, fc300, fc276, fc253, fc231, fc210, fc190, fc171, fc153, fc136, fc120, fc105, fc91, fc78, fc66, fc55, fc45, fc36, fc28, fc21, fc15, fc10, fc6, fc3, fc1, fc0, fs0, in_0_1, in_0_0};

	assign cpa1 = {fc899, fs899, fs898, fs896, fs893, fs889, fs884, fs878, fs871, fs863, fs854, fs844, fs833, fs821, fs808, fs794, fs779, fs763, fs746, fs728, fs709, fs689, fs668, fs646, fs623, fs599, fs574, fs548, fs521, fs493, fs464, fs435, fs406, fs378, fs351, fs325, fs300, fs276, fs253, fs231, fs210, fs190, fs171, fs153, fs136, fs120, fs105, fs91, fs78, fs66, fs55, fs45, fs36, fs28, fs21, fs15, fs10, fs6, fs3, fs1, 1'b0, in_1_0, 1'b0};

	assign res = cpa0 + cpa1;
endmodule
